##
## LEF for PtnCells ;
## created by Innovus v19.11-s128_1 on Sat Sep 10 21:49:25 2022
##

VERSION 5.7 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO DSP
  CLASS BLOCK ;
  SIZE 200.100000 BY 400.520000 ;
  FOREIGN DSP 0.000000 0.000000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN top_N1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 14.5438 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 72.611 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 9.240000 399.820000 9.620000 400.520000 ;
    END
  END top_N1BEG[3]
  PIN top_N1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.0338 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.061 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 7.860000 399.820000 8.240000 400.520000 ;
    END
  END top_N1BEG[2]
  PIN top_N1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.9386 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.585 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 6.480000 399.820000 6.860000 400.520000 ;
    END
  END top_N1BEG[1]
  PIN top_N1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.8 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.892 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 5.100000 399.820000 5.480000 400.520000 ;
    END
  END top_N1BEG[0]
  PIN top_N2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7478 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.631 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 21.660000 399.820000 22.040000 400.520000 ;
    END
  END top_N2BEG[7]
  PIN top_N2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.4146 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.965 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 20.280000 399.820000 20.660000 400.520000 ;
    END
  END top_N2BEG[6]
  PIN top_N2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.4958 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.371 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 18.440000 399.820000 18.820000 400.520000 ;
    END
  END top_N2BEG[5]
  PIN top_N2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7681 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.7325 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 17.060000 399.820000 17.440000 400.520000 ;
    END
  END top_N2BEG[4]
  PIN top_N2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 11.2258 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 56.021 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 15.680000 399.820000 16.060000 400.520000 ;
    END
  END top_N2BEG[3]
  PIN top_N2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.1762 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.773 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 13.840000 399.820000 14.220000 400.520000 ;
    END
  END top_N2BEG[2]
  PIN top_N2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 8.315 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 41.349 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 12.460000 399.820000 12.840000 400.520000 ;
    END
  END top_N2BEG[1]
  PIN top_N2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.0814 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.299 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 11.080000 399.820000 11.460000 400.520000 ;
    END
  END top_N2BEG[0]
  PIN top_N2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2927 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.1845 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 8.8578 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 47.712 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 34.080000 399.820000 34.460000 400.520000 ;
    END
  END top_N2BEGb[7]
  PIN top_N2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.5362 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.455 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 32.240000 399.820000 32.620000 400.520000 ;
    END
  END top_N2BEGb[6]
  PIN top_N2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.917 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.359 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 30.860000 399.820000 31.240000 400.520000 ;
    END
  END top_N2BEGb[5]
  PIN top_N2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.843 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.107 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 29.480000 399.820000 29.860000 400.520000 ;
    END
  END top_N2BEGb[4]
  PIN top_N2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1463 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5705 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.3628 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 29.072 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 27.640000 399.820000 28.020000 400.520000 ;
    END
  END top_N2BEGb[3]
  PIN top_N2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9149 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.4135 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 18.496 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 99.112 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.6678 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.032 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 26.260000 399.820000 26.640000 400.520000 ;
    END
  END top_N2BEGb[2]
  PIN top_N2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7126 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.337 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 24.880000 399.820000 25.260000 400.520000 ;
    END
  END top_N2BEGb[1]
  PIN top_N2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.8414 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.981 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 23.040000 399.820000 23.420000 400.520000 ;
    END
  END top_N2BEGb[0]
  PIN top_N4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 10.9934 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 54.859 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 58.460000 399.820000 58.840000 400.520000 ;
    END
  END top_N4BEG[15]
  PIN top_N4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.1454 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.619 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 56.620000 399.820000 57.000000 400.520000 ;
    END
  END top_N4BEG[14]
  PIN top_N4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.4982 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.383 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 55.240000 399.820000 55.620000 400.520000 ;
    END
  END top_N4BEG[13]
  PIN top_N4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8295 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.9865 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.435 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.12 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 22.8828 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 122.512 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 53.860000 399.820000 54.240000 400.520000 ;
    END
  END top_N4BEG[12]
  PIN top_N4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.4958 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.371 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 52.480000 399.820000 52.860000 400.520000 ;
    END
  END top_N4BEG[11]
  PIN top_N4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.6078 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.931 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 50.640000 399.820000 51.020000 400.520000 ;
    END
  END top_N4BEG[10]
  PIN top_N4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.9869 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.8265 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 49.260000 399.820000 49.640000 400.520000 ;
    END
  END top_N4BEG[9]
  PIN top_N4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7441 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.5595 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.0388 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 27.344 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 47.880000 399.820000 48.260000 400.520000 ;
    END
  END top_N4BEG[8]
  PIN top_N4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1463 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5705 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.9828 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 21.712 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 46.040000 399.820000 46.420000 400.520000 ;
    END
  END top_N4BEG[7]
  PIN top_N4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.479 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.287 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 44.660000 399.820000 45.040000 400.520000 ;
    END
  END top_N4BEG[6]
  PIN top_N4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.115 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.467 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 43.280000 399.820000 43.660000 400.520000 ;
    END
  END top_N4BEG[5]
  PIN top_N4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.1458 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.621 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 41.440000 399.820000 41.820000 400.520000 ;
    END
  END top_N4BEG[4]
  PIN top_N4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.9074 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.429 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 40.060000 399.820000 40.440000 400.520000 ;
    END
  END top_N4BEG[3]
  PIN top_N4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.5434 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.609 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 38.680000 399.820000 39.060000 400.520000 ;
    END
  END top_N4BEG[2]
  PIN top_N4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.9862 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.823 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 36.840000 399.820000 37.220000 400.520000 ;
    END
  END top_N4BEG[1]
  PIN top_N4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.9862 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.823 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 35.460000 399.820000 35.840000 400.520000 ;
    END
  END top_N4BEG[0]
  PIN top_NN4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 7.7167 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 38.4755 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 82.840000 399.820000 83.220000 400.520000 ;
    END
  END top_NN4BEG[15]
  PIN top_NN4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.6702 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 33.243 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 81.460000 399.820000 81.840000 400.520000 ;
    END
  END top_NN4BEG[14]
  PIN top_NN4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.1078 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.313 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 79.620000 399.820000 80.000000 400.520000 ;
    END
  END top_NN4BEG[13]
  PIN top_NN4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.1078 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.313 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 78.240000 399.820000 78.620000 400.520000 ;
    END
  END top_NN4BEG[12]
  PIN top_NN4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.9242 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.513 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 76.860000 399.820000 77.240000 400.520000 ;
    END
  END top_NN4BEG[11]
  PIN top_NN4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.0644 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.096 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 75.020000 399.820000 75.400000 400.520000 ;
    END
  END top_NN4BEG[10]
  PIN top_NN4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.3194 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.489 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 73.640000 399.820000 74.020000 400.520000 ;
    END
  END top_NN4BEG[9]
  PIN top_NN4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.9506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.527 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 72.260000 399.820000 72.640000 400.520000 ;
    END
  END top_NN4BEG[8]
  PIN top_NN4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.2674 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.111 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 70.420000 399.820000 70.800000 400.520000 ;
    END
  END top_NN4BEG[7]
  PIN top_NN4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.9718 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.751 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 69.040000 399.820000 69.420000 400.520000 ;
    END
  END top_NN4BEG[6]
  PIN top_NN4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.0506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.145 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 67.660000 399.820000 68.040000 400.520000 ;
    END
  END top_NN4BEG[5]
  PIN top_NN4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.3838 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.811 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 65.820000 399.820000 66.200000 400.520000 ;
    END
  END top_NN4BEG[4]
  PIN top_NN4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.1465 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.6245 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 64.440000 399.820000 64.820000 400.520000 ;
    END
  END top_NN4BEG[3]
  PIN top_NN4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3853 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.7655 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.6368 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.2 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 63.060000 399.820000 63.440000 400.520000 ;
    END
  END top_NN4BEG[2]
  PIN top_NN4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.2102 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.943 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 61.220000 399.820000 61.600000 400.520000 ;
    END
  END top_NN4BEG[1]
  PIN top_NN4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.4629 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.2065 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 59.840000 399.820000 60.220000 400.520000 ;
    END
  END top_NN4BEG[0]
  PIN top_S1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.5699 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 27.6885 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 17.4594 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 94.048 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.7067 LAYER met3  ;
    ANTENNAMAXAREACAR 43.9464 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 215.215 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 88.820000 399.820000 89.200000 400.520000 ;
    END
  END top_S1END[3]
  PIN top_S1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.2725 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 65.5235 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9117 LAYER met2  ;
    ANTENNAMAXAREACAR 36.6435 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 175.219 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.367145 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 15.4687 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 82.952 LAYER met3  ;
    ANTENNAGATEAREA 1.5477 LAYER met3  ;
    ANTENNAMAXAREACAR 46.6381 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 228.816 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.616411 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 23.2248 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 124.336 LAYER met4  ;
    ANTENNAGATEAREA 1.7067 LAYER met4  ;
    ANTENNAMAXAREACAR 60.2462 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 301.667 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 87.440000 399.820000 87.820000 400.520000 ;
    END
  END top_S1END[2]
  PIN top_S1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 7.0617 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 34.7935 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5937 LAYER met2  ;
    ANTENNAMAXAREACAR 18.5608 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 81.6234 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.532154 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 33.1272 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 177.12 LAYER met3  ;
    ANTENNAGATEAREA 1.5477 LAYER met3  ;
    ANTENNAMAXAREACAR 54.5513 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 271.01 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.616411 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.6698 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 41.376 LAYER met4  ;
    ANTENNAGATEAREA 1.7067 LAYER met4  ;
    ANTENNAMAXAREACAR 59.0452 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 295.253 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 86.060000 399.820000 86.440000 400.520000 ;
    END
  END top_S1END[1]
  PIN top_S1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.0761 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 24.3705 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9117 LAYER met2  ;
    ANTENNAMAXAREACAR 13.8251 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 53.6019 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.411019 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 16.6858 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 89.928 LAYER met3  ;
    ANTENNAGATEAREA 1.3887 LAYER met3  ;
    ANTENNAMAXAREACAR 45.3785 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 221.524 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.577441 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 3.8976 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 21.728 LAYER met4  ;
    ANTENNAGATEAREA 1.7067 LAYER met4  ;
    ANTENNAMAXAREACAR 60.6831 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 306.071 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.47107 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 84.220000 399.820000 84.600000 400.520000 ;
    END
  END top_S1END[0]
  PIN top_S2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 16.8621 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 83.4715 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.0707 LAYER met2  ;
    ANTENNAMAXAREACAR 23.1094 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 108.752 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.502139 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.711 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.592 LAYER met3  ;
    ANTENNAGATEAREA 1.0707 LAYER met3  ;
    ANTENNAMAXAREACAR 24.7074 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 117.711 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.539497 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 42.7932 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 229.632 LAYER met4  ;
    ANTENNAGATEAREA 2.0247 LAYER met4  ;
    ANTENNAMAXAREACAR 99.4453 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 514.78 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 113.200000 399.820000 113.580000 400.520000 ;
    END
  END top_S2MID[7]
  PIN top_S2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.7505 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.4835 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 12.9837 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 46.4182 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.21026 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.255 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 13.5703 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 50.5774 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 76.8354 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 411.2 LAYER met4  ;
    ANTENNAGATEAREA 1.7067 LAYER met4  ;
    ANTENNAMAXAREACAR 118.687 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 623.445 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.952201 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 111.820000 399.820000 112.200000 400.520000 ;
    END
  END top_S2MID[6]
  PIN top_S2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.9759 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.6005 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 10.7723 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 35.0897 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.26202 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.814 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.808 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 12.6448 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 46.1502 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.354037 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 50.8494 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 272.608 LAYER met4  ;
    ANTENNAGATEAREA 1.8657 LAYER met4  ;
    ANTENNAMAXAREACAR 76.2644 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 396.14 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.47107 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 110.440000 399.820000 110.820000 400.520000 ;
    END
  END top_S2MID[5]
  PIN top_S2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 29.1053 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 144.806 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9117 LAYER met2  ;
    ANTENNAMAXAREACAR 50.9362 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 246.132 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.508654 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 11.944 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 64.168 LAYER met3  ;
    ANTENNAGATEAREA 0.9117 LAYER met3  ;
    ANTENNAMAXAREACAR 64.037 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 316.515 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.552528 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 48.2796 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 258.432 LAYER met4  ;
    ANTENNAGATEAREA 1.7067 LAYER met4  ;
    ANTENNAMAXAREACAR 92.3252 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 467.937 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.47107 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 108.600000 399.820000 108.980000 400.520000 ;
    END
  END top_S2MID[4]
  PIN top_S2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.9759 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.6005 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 11.3648 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 38.0527 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.26202 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.471 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 24.312 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 21.6501 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 93.9809 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.354037 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 82.0335 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 438.448 LAYER met4  ;
    ANTENNAGATEAREA 2.0247 LAYER met4  ;
    ANTENNAMAXAREACAR 93.9982 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 478.251 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.637736 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 107.220000 399.820000 107.600000 400.520000 ;
    END
  END top_S2MID[3]
  PIN top_S2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.2705 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.9655 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 9.57902 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 29.1235 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.21026 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.677 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 14.744 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 15.7373 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 63.0412 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 96.5046 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 515.632 LAYER met4  ;
    ANTENNAGATEAREA 1.8657 LAYER met4  ;
    ANTENNAMAXAREACAR 87.5165 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 456.296 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.6587 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 105.840000 399.820000 106.220000 400.520000 ;
    END
  END top_S2MID[2]
  PIN top_S2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.4501 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.9715 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 14.3117 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 52.787 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.26202 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.09 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.28 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 16.8192 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 67.2337 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.354037 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 68.4642 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 367.024 LAYER met4  ;
    ANTENNAGATEAREA 2.0247 LAYER met4  ;
    ANTENNAMAXAREACAR 93.3919 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 483.695 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.967925 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 104.000000 399.820000 104.380000 400.520000 ;
    END
  END top_S2MID[1]
  PIN top_S2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.2171 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.8165 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 11.6085 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 39.5422 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.21026 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.712 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 20.264 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 20.1477 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 86.1583 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 111.914 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 598.272 LAYER met4  ;
    ANTENNAGATEAREA 1.8657 LAYER met4  ;
    ANTENNAMAXAREACAR 98.9662 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 517.505 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 102.620000 399.820000 103.000000 400.520000 ;
    END
  END top_S2MID[0]
  PIN top_S2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 7.1316 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 34.874 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7527 LAYER met2  ;
    ANTENNAMAXAREACAR 17.6274 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 68.9659 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.571064 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 6.227 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 34.144 LAYER met3  ;
    ANTENNAGATEAREA 0.7527 LAYER met3  ;
    ANTENNAMAXAREACAR 25.9003 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 114.328 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.677348 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 12.5226 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 67.728 LAYER met4  ;
    ANTENNAGATEAREA 1.3887 LAYER met4  ;
    ANTENNAMAXAREACAR 39.9363 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 199.855 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 101.240000 399.820000 101.620000 400.520000 ;
    END
  END top_S2END[7]
  PIN top_S2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 10.4828 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 51.919 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7527 LAYER met2  ;
    ANTENNAMAXAREACAR 19.5612 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 79.0184 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.376412 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 14.8017 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 79.408 LAYER met3  ;
    ANTENNAGATEAREA 1.2297 LAYER met3  ;
    ANTENNAMAXAREACAR 31.598 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 143.594 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.574843 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 99.400000 399.820000 99.780000 400.520000 ;
    END
  END top_S2END[6]
  PIN top_S2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.9169 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 34.0795 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5937 LAYER met2  ;
    ANTENNAMAXAREACAR 26.1357 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 123.392 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.532154 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 6.2182 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 33.616 LAYER met3  ;
    ANTENNAGATEAREA 1.0707 LAYER met3  ;
    ANTENNAMAXAREACAR 31.9433 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 154.789 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.612202 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 9.4998 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 51.136 LAYER met4  ;
    ANTENNAGATEAREA 1.2297 LAYER met4  ;
    ANTENNAMAXAREACAR 57.4986 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 295.32 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 98.020000 399.820000 98.400000 400.520000 ;
    END
  END top_S2END[5]
  PIN top_S2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.0303 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.7545 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 15.418 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 58.1171 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.328502 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.09 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.28 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 17.9255 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 72.5638 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.42052 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 32.5818 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 174.24 LAYER met4  ;
    ANTENNAGATEAREA 1.2297 LAYER met4  ;
    ANTENNAMAXAREACAR 46.7671 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 236.327 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.565409 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 96.640000 399.820000 97.020000 400.520000 ;
    END
  END top_S2END[4]
  PIN top_S2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0276 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.977 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.884 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 15.848 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 21.6966 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 116.656 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3887 LAYER met4  ;
    ANTENNAMAXAREACAR 72.6426 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 361.758 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.663897 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 95.260000 399.820000 95.640000 400.520000 ;
    END
  END top_S2END[3]
  PIN top_S2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.2457 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 25.9595 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 18.0529 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 71.7644 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.21026 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.447 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 24.184 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 28.283 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 127.398 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 22.5573 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 121.712 LAYER met4  ;
    ANTENNAGATEAREA 1.3887 LAYER met4  ;
    ANTENNAMAXAREACAR 65.9542 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 341.5 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.47107 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 93.420000 399.820000 93.800000 400.520000 ;
    END
  END top_S2END[2]
  PIN top_S2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3853 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.7655 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 20.4634 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 109.6 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9117 LAYER met3  ;
    ANTENNAMAXAREACAR 49.6125 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 248.404 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.411019 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 23.2248 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 124.336 LAYER met4  ;
    ANTENNAGATEAREA 1.3887 LAYER met4  ;
    ANTENNAMAXAREACAR 66.3366 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 337.938 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.632495 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 92.040000 399.820000 92.420000 400.520000 ;
    END
  END top_S2END[1]
  PIN top_S2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.1229 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 24.7555 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9117 LAYER met2  ;
    ANTENNAMAXAREACAR 27.2313 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 128.1 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.650163 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.2509 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAGATEAREA 0.9117 LAYER met3  ;
    ANTENNAMAXAREACAR 27.5065 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 130.083 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.694037 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 37.2048 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 198.896 LAYER met4  ;
    ANTENNAGATEAREA 1.3887 LAYER met4  ;
    ANTENNAMAXAREACAR 54.2976 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 273.307 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.694037 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 90.660000 399.820000 91.040000 400.520000 ;
    END
  END top_S2END[0]
  PIN top_S4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1711 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.6945 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.472 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 34.984 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.3041 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 114.239 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 610.688 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.5006 LAYER met4  ;
    ANTENNAMAXAREACAR 107.831 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 571.309 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.19033 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 138.040000 399.820000 138.420000 400.520000 ;
    END
  END top_S4END[15]
  PIN top_S4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9435 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.5565 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.3041 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 115.095 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 614.304 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.5006 LAYER met4  ;
    ANTENNAMAXAREACAR 89.8684 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 458.843 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 136.200000 399.820000 136.580000 400.520000 ;
    END
  END top_S4END[14]
  PIN top_S4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9149 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.4135 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.366 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.752 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.3041 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 115.927 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 619.216 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.5006 LAYER met4  ;
    ANTENNAMAXAREACAR 110.912 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 591.058 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.872265 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 134.820000 399.820000 135.200000 400.520000 ;
    END
  END top_S4END[13]
  PIN top_S4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8581 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.1295 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.435 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.12 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.3041 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 111.44 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 594.816 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.5006 LAYER met4  ;
    ANTENNAMAXAREACAR 81.0144 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 412.158 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.31489 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 133.440000 399.820000 133.820000 400.520000 ;
    END
  END top_S4END[12]
  PIN top_S4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7479 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.5785 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.676 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.072 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.3041 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 112.379 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 599.824 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.5006 LAYER met4  ;
    ANTENNAMAXAREACAR 86.0248 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 444.053 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.491796 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 131.600000 399.820000 131.980000 400.520000 ;
    END
  END top_S4END[11]
  PIN top_S4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0647 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.1625 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.918 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.696 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.8694 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 114.374 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 611.408 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.0659 LAYER met4  ;
    ANTENNAMAXAREACAR 124.661 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 659.698 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.591883 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 130.220000 399.820000 130.600000 400.520000 ;
    END
  END top_S4END[10]
  PIN top_S4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6835 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.2565 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.9008 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 32.408 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 90.8718 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 485.12 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6312 LAYER met4  ;
    ANTENNAMAXAREACAR 159.065 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 826.719 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.38832 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 128.840000 399.820000 129.220000 400.520000 ;
    END
  END top_S4END[9]
  PIN top_S4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.2717 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 26.1975 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.135 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.52 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 101.581 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 544.112 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6312 LAYER met4  ;
    ANTENNAMAXAREACAR 181.76 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 965.56 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 127.000000 399.820000 127.380000 400.520000 ;
    END
  END top_S4END[8]
  PIN top_S4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.1393 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 25.4275 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 15.9156 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 61.233 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.21026 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 16.8357 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 67.2142 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 91.5561 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 490.176 LAYER met4  ;
    ANTENNAGATEAREA 1.2297 LAYER met4  ;
    ANTENNAMAXAREACAR 128.281 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 667.404 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.32956 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 125.620000 399.820000 126.000000 400.520000 ;
    END
  END top_S4END[7]
  PIN top_S4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.8965 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.2135 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 10.7562 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 35.4359 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.21026 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.745 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.44 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 12.47 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 45.6499 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 90.4254 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 483.68 LAYER met4  ;
    ANTENNAGATEAREA 1.2297 LAYER met4  ;
    ANTENNAMAXAREACAR 131.932 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 685.574 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.07799 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 124.240000 399.820000 124.620000 400.520000 ;
    END
  END top_S4END[6]
  PIN top_S4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.4561 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 22.0115 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 14.4587 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 53.7934 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.21026 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.368 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 29.096 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 26.8075 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 120.727 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 86.1378 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 459.872 LAYER met4  ;
    ANTENNAGATEAREA 1.2297 LAYER met4  ;
    ANTENNAMAXAREACAR 106.43 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 547.281 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.706918 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 122.400000 399.820000 122.780000 400.520000 ;
    END
  END top_S4END[5]
  PIN top_S4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.4761 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.1015 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 9.02991 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 26.378 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.26202 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.09 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.28 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 11.5374 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 40.8247 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.354037 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 89.5506 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 478.544 LAYER met4  ;
    ANTENNAGATEAREA 1.2297 LAYER met4  ;
    ANTENNAMAXAREACAR 117.936 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 610.516 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.682809 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 121.020000 399.820000 121.400000 400.520000 ;
    END
  END top_S4END[4]
  PIN top_S4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.1923 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.6925 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 9.84357 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 30.7177 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.21026 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.2509 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 10.4207 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 34.8769 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 23.8056 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 127.904 LAYER met4  ;
    ANTENNAGATEAREA 1.2297 LAYER met4  ;
    ANTENNAMAXAREACAR 55.712 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 278.903 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 119.640000 399.820000 120.020000 400.520000 ;
    END
  END top_S4END[3]
  PIN top_S4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.6079 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.6525 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 10.0922 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 31.8449 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.21026 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.264 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 23.208 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 19.9013 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 85.2335 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 28.5558 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 152.768 LAYER met4  ;
    ANTENNAGATEAREA 1.2297 LAYER met4  ;
    ANTENNAMAXAREACAR 67.0869 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 342.364 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.682809 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 117.800000 399.820000 118.180000 400.520000 ;
    END
  END top_S4END[2]
  PIN top_S4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1463 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5705 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.642 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.224 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 33.9348 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 181.456 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2297 LAYER met4  ;
    ANTENNAMAXAREACAR 72.946 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 367.826 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.74888 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 116.420000 399.820000 116.800000 400.520000 ;
    END
  END top_S4END[1]
  PIN top_S4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.0673 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.0675 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 11.1491 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 37.4005 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.21026 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.298 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 18.056 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 18.7359 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 78.9372 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 19.7076 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 106.048 LAYER met4  ;
    ANTENNAGATEAREA 1.2297 LAYER met4  ;
    ANTENNAMAXAREACAR 72.1516 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 368.698 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 115.040000 399.820000 115.420000 400.520000 ;
    END
  END top_S4END[0]
  PIN top_SS4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9397 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.5375 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.85 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 21 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.3041 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 112.697 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 601.52 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.5006 LAYER met4  ;
    ANTENNAMAXAREACAR 88.0606 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 448.165 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.491796 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 162.420000 399.820000 162.800000 400.520000 ;
    END
  END top_SS4END[15]
  PIN top_SS4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9645 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.6615 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.574 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 19.528 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.3041 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 111.082 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 593.376 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.5006 LAYER met4  ;
    ANTENNAMAXAREACAR 82.7387 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 418.257 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 160.580000 399.820000 160.960000 400.520000 ;
    END
  END top_SS4END[14]
  PIN top_SS4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7689 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.6835 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.01 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 32.52 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.7388 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 116.62 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 622.912 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.9353 LAYER met4  ;
    ANTENNAMAXAREACAR 67.5743 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 351.95 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 159.200000 399.820000 159.580000 400.520000 ;
    END
  END top_SS4END[13]
  PIN top_SS4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.2245 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 20.9615 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.918 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.696 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 101.934 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 544.112 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6312 LAYER met4  ;
    ANTENNAMAXAREACAR 188.482 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 995.773 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 157.820000 399.820000 158.200000 400.520000 ;
    END
  END top_SS4END[12]
  PIN top_SS4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1463 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5705 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.129 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 54.488 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.7388 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 118.125 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 630.464 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.9353 LAYER met4  ;
    ANTENNAMAXAREACAR 67.3616 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 356.381 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 155.980000 399.820000 156.360000 400.520000 ;
    END
  END top_SS4END[11]
  PIN top_SS4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8295 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.9865 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.676 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.072 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.3041 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 120.208 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 642.048 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.5006 LAYER met4  ;
    ANTENNAMAXAREACAR 96.8035 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 495.762 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.872265 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 154.600000 399.820000 154.980000 400.520000 ;
    END
  END top_SS4END[10]
  PIN top_SS4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1463 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5705 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.3041 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 117.137 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 625.2 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.5006 LAYER met4  ;
    ANTENNAMAXAREACAR 90.0459 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 467.926 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.491796 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 153.220000 399.820000 153.600000 400.520000 ;
    END
  END top_SS4END[9]
  PIN top_SS4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3419 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.5485 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.022 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 16.584 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.8694 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 110.398 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 589.728 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.0659 LAYER met4  ;
    ANTENNAMAXAREACAR 155.043 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 816.616 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.872265 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 151.380000 399.820000 151.760000 400.520000 ;
    END
  END top_SS4END[8]
  PIN top_SS4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.2171 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.8165 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 11.6085 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 39.5422 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.21026 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.195 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 22.84 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 21.2588 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 92.0842 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 85.7718 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 457.92 LAYER met4  ;
    ANTENNAGATEAREA 0.7527 LAYER met4  ;
    ANTENNAMAXAREACAR 135.211 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 700.454 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.574843 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 150.000000 399.820000 150.380000 400.520000 ;
    END
  END top_SS4END[7]
  PIN top_SS4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.8321 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.8915 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 10.608 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 34.6952 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.21026 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.538 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.336 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 11.8456 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 42.3694 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 83.0898 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 443.616 LAYER met4  ;
    ANTENNAGATEAREA 0.9117 LAYER met4  ;
    ANTENNAMAXAREACAR 169.064 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 885.957 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.6587 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 148.620000 399.820000 149.000000 400.520000 ;
    END
  END top_SS4END[6]
  PIN top_SS4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.4979 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.0925 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 13.7509 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 49.7113 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.26202 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.78 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.96 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 17.8456 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 72.6236 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.354037 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 72.3966 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 387.056 LAYER met4  ;
    ANTENNAGATEAREA 0.9117 LAYER met4  ;
    ANTENNAMAXAREACAR 165.529 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 875.48 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.07799 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 146.780000 399.820000 147.160000 400.520000 ;
    END
  END top_SS4END[5]
  PIN top_SS4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.1069 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.2655 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 8.93973 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 26.3538 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.21026 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.255 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 9.52634 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 30.513 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 110.502 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 592.16 LAYER met4  ;
    ANTENNAGATEAREA 0.9117 LAYER met4  ;
    ANTENNAMAXAREACAR 143.324 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 757.487 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.32956 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 145.400000 399.820000 145.780000 400.520000 ;
    END
  END top_SS4END[4]
  PIN top_SS4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1463 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5705 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 9.8068 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 53.24 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 34.2742 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 162.557 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.394295 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 13.3188 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 71.504 LAYER met4  ;
    ANTENNAGATEAREA 0.7527 LAYER met4  ;
    ANTENNAMAXAREACAR 60.9145 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 305.813 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.574843 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 144.020000 399.820000 144.400000 400.520000 ;
    END
  END top_SS4END[3]
  PIN top_SS4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.2325 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 20.7655 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 16.9618 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 65.766 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.26202 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.2509 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 17.539 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 69.9252 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.354037 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 20.8524 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 112.624 LAYER met4  ;
    ANTENNAGATEAREA 0.9117 LAYER met4  ;
    ANTENNAMAXAREACAR 97.9701 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 516.107 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.32956 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 142.640000 399.820000 143.020000 400.520000 ;
    END
  END top_SS4END[2]
  PIN top_SS4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.6781 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.9935 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 19.2206 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 77.2153 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.26202 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.987 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.064 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 23.7916 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 102.667 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.354037 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 23.2314 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 125.312 LAYER met4  ;
    ANTENNAGATEAREA 0.9117 LAYER met4  ;
    ANTENNAMAXAREACAR 93.0584 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 493.273 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.07799 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 140.800000 399.820000 141.180000 400.520000 ;
    END
  END top_SS4END[1]
  PIN top_SS4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.3423 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.4325 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 13.4663 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 48.5599 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.26202 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.9629 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 16.264 LAYER met3  ;
    ANTENNAGATEAREA 0.5937 LAYER met3  ;
    ANTENNAMAXAREACAR 18.4569 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 75.9542 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.642217 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 19.0464 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 102.992 LAYER met4  ;
    ANTENNAGATEAREA 0.9117 LAYER met4  ;
    ANTENNAMAXAREACAR 67.9068 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 350.973 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 139.420000 399.820000 139.800000 400.520000 ;
    END
  END top_SS4END[0]
  PIN top_E1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.5064 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 18.696 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 280.800000 200.100000 281.180000 ;
    END
  END top_E1BEG[3]
  PIN top_E1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 279.580000 200.100000 279.960000 ;
    END
  END top_E1BEG[2]
  PIN top_E1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.1264 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.336 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 277.750000 200.100000 278.130000 ;
    END
  END top_E1BEG[1]
  PIN top_E1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 276.530000 200.100000 276.910000 ;
    END
  END top_E1BEG[0]
  PIN top_E2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.8614 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 15.256 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 293.000000 200.100000 293.380000 ;
    END
  END top_E2BEG[7]
  PIN top_E2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 291.170000 200.100000 291.550000 ;
    END
  END top_E2BEG[6]
  PIN top_E2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 289.950000 200.100000 290.330000 ;
    END
  END top_E2BEG[5]
  PIN top_E2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 288.120000 200.100000 288.500000 ;
    END
  END top_E2BEG[4]
  PIN top_E2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.8164 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 15.016 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 286.900000 200.100000 287.280000 ;
    END
  END top_E2BEG[3]
  PIN top_E2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 285.070000 200.100000 285.450000 ;
    END
  END top_E2BEG[2]
  PIN top_E2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.4364 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.656 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 283.850000 200.100000 284.230000 ;
    END
  END top_E2BEG[1]
  PIN top_E2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 282.020000 200.100000 282.400000 ;
    END
  END top_E2BEG[0]
  PIN top_E2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 304.590000 200.100000 304.970000 ;
    END
  END top_E2BEGb[7]
  PIN top_E2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.8844 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.712 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 303.370000 200.100000 303.750000 ;
    END
  END top_E2BEGb[6]
  PIN top_E2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.8934 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.76 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 301.540000 200.100000 301.920000 ;
    END
  END top_E2BEGb[5]
  PIN top_E2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.2984 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.92 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 300.320000 200.100000 300.700000 ;
    END
  END top_E2BEGb[4]
  PIN top_E2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 298.490000 200.100000 298.870000 ;
    END
  END top_E2BEGb[3]
  PIN top_E2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 297.270000 200.100000 297.650000 ;
    END
  END top_E2BEGb[2]
  PIN top_E2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.9884 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.28 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 295.440000 200.100000 295.820000 ;
    END
  END top_E2BEGb[1]
  PIN top_E2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.1604 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.184 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 294.220000 200.100000 294.600000 ;
    END
  END top_E2BEGb[0]
  PIN top_EE4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 328.380000 200.100000 328.760000 ;
    END
  END top_EE4BEG[15]
  PIN top_EE4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.4364 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.656 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 327.160000 200.100000 327.540000 ;
    END
  END top_EE4BEG[14]
  PIN top_EE4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 325.330000 200.100000 325.710000 ;
    END
  END top_EE4BEG[13]
  PIN top_EE4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.7124 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.128 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 324.110000 200.100000 324.490000 ;
    END
  END top_EE4BEG[12]
  PIN top_EE4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.4364 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.656 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 322.280000 200.100000 322.660000 ;
    END
  END top_EE4BEG[11]
  PIN top_EE4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 321.060000 200.100000 321.440000 ;
    END
  END top_EE4BEG[10]
  PIN top_EE4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.3344 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 23.112 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 319.230000 200.100000 319.610000 ;
    END
  END top_EE4BEG[9]
  PIN top_EE4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 318.010000 200.100000 318.390000 ;
    END
  END top_EE4BEG[8]
  PIN top_EE4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.8504 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.864 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 316.790000 200.100000 317.170000 ;
    END
  END top_EE4BEG[7]
  PIN top_EE4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 314.960000 200.100000 315.340000 ;
    END
  END top_EE4BEG[6]
  PIN top_EE4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.2644 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 12.072 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 313.740000 200.100000 314.120000 ;
    END
  END top_EE4BEG[5]
  PIN top_EE4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 311.910000 200.100000 312.290000 ;
    END
  END top_EE4BEG[4]
  PIN top_EE4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.7124 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.128 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 310.690000 200.100000 311.070000 ;
    END
  END top_EE4BEG[3]
  PIN top_EE4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.5744 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.392 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 308.860000 200.100000 309.240000 ;
    END
  END top_EE4BEG[2]
  PIN top_EE4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.4364 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.656 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 307.640000 200.100000 308.020000 ;
    END
  END top_EE4BEG[1]
  PIN top_EE4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 305.810000 200.100000 306.190000 ;
    END
  END top_EE4BEG[0]
  PIN top_E6BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.6084 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.24 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 346.070000 200.100000 346.450000 ;
    END
  END top_E6BEG[11]
  PIN top_E6BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 344.850000 200.100000 345.230000 ;
    END
  END top_E6BEG[10]
  PIN top_E6BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.7124 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.128 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 343.630000 200.100000 344.010000 ;
    END
  END top_E6BEG[9]
  PIN top_E6BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 341.800000 200.100000 342.180000 ;
    END
  END top_E6BEG[8]
  PIN top_E6BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.6444 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 19.432 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 340.580000 200.100000 340.960000 ;
    END
  END top_E6BEG[7]
  PIN top_E6BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.1604 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.184 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 338.750000 200.100000 339.130000 ;
    END
  END top_E6BEG[6]
  PIN top_E6BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 6.1284 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 32.68 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 337.530000 200.100000 337.910000 ;
    END
  END top_E6BEG[5]
  PIN top_E6BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.4724 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 23.848 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 335.700000 200.100000 336.080000 ;
    END
  END top_E6BEG[4]
  PIN top_E6BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 334.480000 200.100000 334.860000 ;
    END
  END top_E6BEG[3]
  PIN top_E6BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 332.650000 200.100000 333.030000 ;
    END
  END top_E6BEG[2]
  PIN top_E6BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 331.430000 200.100000 331.810000 ;
    END
  END top_E6BEG[1]
  PIN top_E6BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.7464 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.976 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 330.210000 200.100000 330.590000 ;
    END
  END top_E6BEG[0]
  PIN top_E1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 31.2049 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 167.344 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.7067 LAYER met3  ;
    ANTENNAMAXAREACAR 57.0044 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 283.144 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.59828 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 10.5336 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 57.12 LAYER met4  ;
    ANTENNAGATEAREA 2.1837 LAYER met4  ;
    ANTENNAMAXAREACAR 61.8282 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 309.302 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.07799 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 280.800000 0.700000 281.180000 ;
    END
  END top_E1END[3]
  PIN top_E1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.435 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 39.64 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.318 LAYER met3  ;
    ANTENNAMAXAREACAR 42.1167 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 210.008 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.574843 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 22.8012 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 123.488 LAYER met4  ;
    ANTENNAGATEAREA 2.1837 LAYER met4  ;
    ANTENNAMAXAREACAR 52.5582 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 266.558 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.02553 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 279.580000 0.700000 279.960000 ;
    END
  END top_E1END[2]
  PIN top_E1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 20.2821 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 108.632 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.8657 LAYER met3  ;
    ANTENNAMAXAREACAR 34.8926 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 172.798 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.490625 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 277.750000 0.700000 278.130000 ;
    END
  END top_E1END[1]
  PIN top_E1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.7296 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 25.216 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 20.4864 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 110.672 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.8657 LAYER met4  ;
    ANTENNAMAXAREACAR 75.3824 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 389.716 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.967925 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 276.530000 0.700000 276.910000 ;
    END
  END top_E1END[0]
  PIN top_E2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 26.5114 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 141.856 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 6.0102 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 36.288 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8325 LAYER met4  ;
    ANTENNAMAXAREACAR 51.7239 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 272.121 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.72264 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 293.000000 0.700000 293.380000 ;
    END
  END top_E2MID[7]
  PIN top_E2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 29.239 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 156.408 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 13.1361 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 71.936 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6735 LAYER met4  ;
    ANTENNAMAXAREACAR 43.3317 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 219 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 291.170000 0.700000 291.550000 ;
    END
  END top_E2MID[6]
  PIN top_E2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.4981 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 18.528 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.5828 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.912 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8325 LAYER met4  ;
    ANTENNAMAXAREACAR 85.7157 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 442.87 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.680543 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 289.950000 0.700000 290.330000 ;
    END
  END top_E2MID[5]
  PIN top_E2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 20.5486 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 109.584 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.9488 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 10.864 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6735 LAYER met4  ;
    ANTENNAMAXAREACAR 69.8808 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 357.827 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.885806 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 288.120000 0.700000 288.500000 ;
    END
  END top_E2MID[4]
  PIN top_E2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.6596 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 14.176 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 3.2844 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 18.928 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8325 LAYER met4  ;
    ANTENNAMAXAREACAR 76.7345 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 397.579 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.716352 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 286.900000 0.700000 287.280000 ;
    END
  END top_E2MID[3]
  PIN top_E2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8316 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 25.76 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.7354 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 16 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6735 LAYER met4  ;
    ANTENNAMAXAREACAR 22.9949 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 114.05 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.634234 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 285.070000 0.700000 285.450000 ;
    END
  END top_E2MID[2]
  PIN top_E2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.9476 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 31.712 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 6.6972 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 37.6 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8325 LAYER met4  ;
    ANTENNAMAXAREACAR 77.1279 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 388.774 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.921633 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 283.850000 0.700000 284.230000 ;
    END
  END top_E2MID[1]
  PIN top_E2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.6124 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 78.376 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.477 LAYER met3  ;
    ANTENNAMAXAREACAR 70.2537 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 351.932 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.716352 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 4.437 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 26.016 LAYER met4  ;
    ANTENNAGATEAREA 0.6735 LAYER met4  ;
    ANTENNAMAXAREACAR 76.8417 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 390.56 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.716352 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 282.020000 0.700000 282.400000 ;
    END
  END top_E2MID[0]
  PIN top_E2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 35.571 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 190.648 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2297 LAYER met3  ;
    ANTENNAMAXAREACAR 54.0531 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 261.752 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.716352 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 304.590000 0.700000 304.970000 ;
    END
  END top_E2END[7]
  PIN top_E2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.4766 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 13.2 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 29.0166 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 155.696 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3887 LAYER met4  ;
    ANTENNAMAXAREACAR 54.6735 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 283.319 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04264 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 303.370000 0.700000 303.750000 ;
    END
  END top_E2END[6]
  PIN top_E2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3887 LAYER met3  ;
    ANTENNAMAXAREACAR 62.1938 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 302.076 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.635093 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 301.540000 0.700000 301.920000 ;
    END
  END top_E2END[5]
  PIN top_E2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.4766 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 13.2 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 14.3298 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 76.896 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2297 LAYER met4  ;
    ANTENNAMAXAREACAR 28.591 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 128.79 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.529836 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 300.320000 0.700000 300.700000 ;
    END
  END top_E2END[4]
  PIN top_E2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 12.9582 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 69.576 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.7067 LAYER met3  ;
    ANTENNAMAXAREACAR 33.9988 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 162.917 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.488217 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 298.490000 0.700000 298.870000 ;
    END
  END top_E2END[3]
  PIN top_E2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 23.9631 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 128.264 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.5477 LAYER met3  ;
    ANTENNAMAXAREACAR 44.2374 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 218.732 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.574843 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 297.270000 0.700000 297.650000 ;
    END
  END top_E2END[2]
  PIN top_E2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 20.476 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 109.672 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9117 LAYER met3  ;
    ANTENNAMAXAREACAR 44.9038 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 213.557 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.596402 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.8508 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 5.008 LAYER met4  ;
    ANTENNAGATEAREA 1.0707 LAYER met4  ;
    ANTENNAMAXAREACAR 45.6984 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 218.235 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 295.440000 0.700000 295.820000 ;
    END
  END top_E2END[1]
  PIN top_E2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0736 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 16.384 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 59.6673 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 319.632 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.0707 LAYER met4  ;
    ANTENNAMAXAREACAR 85.8768 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 451.509 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.884067 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 294.220000 0.700000 294.600000 ;
    END
  END top_E2END[0]
  PIN top_EE4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.09 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.265 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 14.432 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 48.6662 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 262.265 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 328.380000 0.700000 328.760000 ;
    END
  END top_EE4END[15]
  PIN top_EE4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 48.7006 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 259.728 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.3356 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.064 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 34.0422 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 180.672 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 327.160000 0.700000 327.540000 ;
    END
  END top_EE4END[14]
  PIN top_EE4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 49.7794 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 265.952 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.6166 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 14.896 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 34.5934 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 185.293 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 325.330000 0.700000 325.710000 ;
    END
  END top_EE4END[13]
  PIN top_EE4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 49.0024 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 261.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.3052 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 14.176 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 38.2204 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 203.232 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 324.110000 0.700000 324.490000 ;
    END
  END top_EE4END[12]
  PIN top_EE4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 50.0386 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 266.864 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.9696 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 6.112 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 24.7659 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 131.796 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 322.280000 0.700000 322.660000 ;
    END
  END top_EE4END[11]
  PIN top_EE4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 36.9544 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 197.552 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.9696 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 6.112 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 20.9043 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 113.308 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 321.060000 0.700000 321.440000 ;
    END
  END top_EE4END[10]
  PIN top_EE4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.2164 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 17.616 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 12.3942 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 67.984 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 97.1903 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 515.98 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 319.230000 0.700000 319.610000 ;
    END
  END top_EE4END[9]
  PIN top_EE4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 43.426 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 232.072 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.6614 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 10.272 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 28.0209 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 150.025 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 318.010000 0.700000 318.390000 ;
    END
  END top_EE4END[8]
  PIN top_EE4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 32.6764 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 174.736 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.3356 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.064 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 37.3659 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 197.45 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 316.790000 0.700000 317.170000 ;
    END
  END top_EE4END[7]
  PIN top_EE4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 50.5306 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 269.488 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.4336 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 13.92 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 37.2361 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 194.662 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 314.960000 0.700000 315.340000 ;
    END
  END top_EE4END[6]
  PIN top_EE4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 52.7764 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 281.936 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.1864 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 13.072 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 30.712 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 166.57 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 313.740000 0.700000 314.120000 ;
    END
  END top_EE4END[5]
  PIN top_EE4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 41.176 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 220.072 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.2954 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.32 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 36.6112 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 192.087 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 311.910000 0.700000 312.290000 ;
    END
  END top_EE4END[4]
  PIN top_EE4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 9.9994 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 53.792 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 34.5466 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 162.547 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.446055 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.4848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 3.056 LAYER met4  ;
    ANTENNAGATEAREA 0.7527 LAYER met4  ;
    ANTENNAMAXAREACAR 61.1658 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 311.257 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.716352 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 310.690000 0.700000 311.070000 ;
    END
  END top_EE4END[3]
  PIN top_EE4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 45.9793 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 245.68 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5937 LAYER met3  ;
    ANTENNAMAXAREACAR 92.3453 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 469.666 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.642217 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 9.8517 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 53.008 LAYER met4  ;
    ANTENNAGATEAREA 0.9117 LAYER met4  ;
    ANTENNAMAXAREACAR 103.151 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 527.808 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 308.860000 0.700000 309.240000 ;
    END
  END top_EE4END[2]
  PIN top_EE4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 17.9041 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 96.416 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7527 LAYER met3  ;
    ANTENNAMAXAREACAR 52.8301 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 266.465 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.879557 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 3.0468 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 16.72 LAYER met4  ;
    ANTENNAGATEAREA 0.9117 LAYER met4  ;
    ANTENNAMAXAREACAR 56.1719 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 284.804 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.879557 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 307.640000 0.700000 308.020000 ;
    END
  END top_EE4END[1]
  PIN top_EE4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.0282 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 74.8 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 11.1774 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 61.024 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9117 LAYER met4  ;
    ANTENNAMAXAREACAR 46.7179 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 233.551 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 305.810000 0.700000 306.190000 ;
    END
  END top_EE4END[0]
  PIN top_E6END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.4786 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 18.544 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 19.7928 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 108.384 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6312 LAYER met4  ;
    ANTENNAMAXAREACAR 80.6642 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 416.007 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.846577 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 346.070000 0.700000 346.450000 ;
    END
  END top_E6END[11]
  PIN top_E6END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 38.602 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 206.344 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.9696 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 6.112 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 15.1593 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 84.5394 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 344.850000 0.700000 345.230000 ;
    END
  END top_E6END[10]
  PIN top_E6END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 51.3196 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 273.696 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.9696 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 6.112 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 21.685 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 116.626 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 343.630000 0.700000 344.010000 ;
    END
  END top_E6END[9]
  PIN top_E6END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.6412 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 79.032 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 84.1776 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 446.621 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.46514 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 341.800000 0.700000 342.180000 ;
    END
  END top_E6END[8]
  PIN top_E6END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3534 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.68 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 3.9618 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 21.6 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 26.6626 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 141.517 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 340.580000 0.700000 340.960000 ;
    END
  END top_E6END[7]
  PIN top_E6END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 46.4476 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 247.712 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.9696 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 6.112 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 30.17 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 153.435 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 338.750000 0.700000 339.130000 ;
    END
  END top_E6END[6]
  PIN top_E6END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 48.5176 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 258.752 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.7016 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 10.016 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 20.5099 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 111.608 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 337.530000 0.700000 337.910000 ;
    END
  END top_E6END[5]
  PIN top_E6END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 51.3196 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 273.696 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.7016 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 10.016 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 28.6738 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 153.598 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 335.700000 0.700000 336.080000 ;
    END
  END top_E6END[4]
  PIN top_E6END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 48.028 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 256.616 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.9696 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 6.112 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 33.6952 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 173.939 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 334.480000 0.700000 334.860000 ;
    END
  END top_E6END[3]
  PIN top_E6END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.6664 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 212.016 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.3356 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.064 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 19.885 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 107.471 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 332.650000 0.700000 333.030000 ;
    END
  END top_E6END[2]
  PIN top_E6END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 7.2039 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 39.352 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.3427 LAYER met3  ;
    ANTENNAMAXAREACAR 36.754 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 174.155 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.967925 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 331.430000 0.700000 331.810000 ;
    END
  END top_E6END[1]
  PIN top_E6END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.7292 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 25.688 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.3427 LAYER met3  ;
    ANTENNAMAXAREACAR 70.2879 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 343.719 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.634242 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 330.210000 0.700000 330.590000 ;
    END
  END top_E6END[0]
  PIN top_W1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 209.430000 0.700000 209.810000 ;
    END
  END top_W1BEG[3]
  PIN top_W1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.9204 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 20.904 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 207.600000 0.700000 207.980000 ;
    END
  END top_W1BEG[2]
  PIN top_W1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 206.380000 0.700000 206.760000 ;
    END
  END top_W1BEG[1]
  PIN top_W1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.6444 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 19.432 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 205.160000 0.700000 205.540000 ;
    END
  END top_W1BEG[0]
  PIN top_W2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 38.7882 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 207.816 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 221.020000 0.700000 221.400000 ;
    END
  END top_W2BEG[7]
  PIN top_W2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 219.800000 0.700000 220.180000 ;
    END
  END top_W2BEG[6]
  PIN top_W2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.4724 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 23.848 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 217.970000 0.700000 218.350000 ;
    END
  END top_W2BEG[5]
  PIN top_W2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 216.750000 0.700000 217.130000 ;
    END
  END top_W2BEG[4]
  PIN top_W2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 14.9094 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 79.512 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 215.530000 0.700000 215.910000 ;
    END
  END top_W2BEG[3]
  PIN top_W2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 213.700000 0.700000 214.080000 ;
    END
  END top_W2BEG[2]
  PIN top_W2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.6084 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.24 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 212.480000 0.700000 212.860000 ;
    END
  END top_W2BEG[1]
  PIN top_W2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 12.8874 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 68.728 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 210.650000 0.700000 211.030000 ;
    END
  END top_W2BEG[0]
  PIN top_W2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 35.0622 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 187.944 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 233.220000 0.700000 233.600000 ;
    END
  END top_W2BEGb[7]
  PIN top_W2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 28.2924 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 150.888 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 231.390000 0.700000 231.770000 ;
    END
  END top_W2BEGb[6]
  PIN top_W2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 230.170000 0.700000 230.550000 ;
    END
  END top_W2BEGb[5]
  PIN top_W2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.2984 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.92 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 228.950000 0.700000 229.330000 ;
    END
  END top_W2BEGb[4]
  PIN top_W2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 11.3244 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 60.392 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 227.120000 0.700000 227.500000 ;
    END
  END top_W2BEGb[3]
  PIN top_W2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 17.2278 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 92.352 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 225.900000 0.700000 226.280000 ;
    END
  END top_W2BEGb[2]
  PIN top_W2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.1296 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 166.016 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.6678 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.032 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 224.070000 0.700000 224.450000 ;
    END
  END top_W2BEGb[1]
  PIN top_W2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 222.850000 0.700000 223.230000 ;
    END
  END top_W2BEGb[0]
  PIN top_WW4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.8844 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.712 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 257.010000 0.700000 257.390000 ;
    END
  END top_WW4BEG[15]
  PIN top_WW4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 255.180000 0.700000 255.560000 ;
    END
  END top_WW4BEG[14]
  PIN top_WW4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.9544 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 15.752 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 253.960000 0.700000 254.340000 ;
    END
  END top_WW4BEG[13]
  PIN top_WW4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 252.740000 0.700000 253.120000 ;
    END
  END top_WW4BEG[12]
  PIN top_WW4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 250.910000 0.700000 251.290000 ;
    END
  END top_WW4BEG[11]
  PIN top_WW4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 249.690000 0.700000 250.070000 ;
    END
  END top_WW4BEG[10]
  PIN top_WW4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.3684 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 17.96 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 247.860000 0.700000 248.240000 ;
    END
  END top_WW4BEG[9]
  PIN top_WW4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 246.640000 0.700000 247.020000 ;
    END
  END top_WW4BEG[8]
  PIN top_WW4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 244.810000 0.700000 245.190000 ;
    END
  END top_WW4BEG[7]
  PIN top_WW4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.6084 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.24 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 243.590000 0.700000 243.970000 ;
    END
  END top_WW4BEG[6]
  PIN top_WW4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.0224 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.448 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 242.370000 0.700000 242.750000 ;
    END
  END top_WW4BEG[5]
  PIN top_WW4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.5404 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 13.544 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 240.540000 0.700000 240.920000 ;
    END
  END top_WW4BEG[4]
  PIN top_WW4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 239.320000 0.700000 239.700000 ;
    END
  END top_WW4BEG[3]
  PIN top_WW4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.9544 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 15.752 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 237.490000 0.700000 237.870000 ;
    END
  END top_WW4BEG[2]
  PIN top_WW4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 236.270000 0.700000 236.650000 ;
    END
  END top_WW4BEG[1]
  PIN top_WW4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.1604 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.184 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 234.440000 0.700000 234.820000 ;
    END
  END top_WW4BEG[0]
  PIN top_W6BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.5864 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.312 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 274.700000 0.700000 275.080000 ;
    END
  END top_W6BEG[11]
  PIN top_W6BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 273.480000 0.700000 273.860000 ;
    END
  END top_W6BEG[10]
  PIN top_W6BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.2504 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.664 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 271.650000 0.700000 272.030000 ;
    END
  END top_W6BEG[9]
  PIN top_W6BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 270.430000 0.700000 270.810000 ;
    END
  END top_W6BEG[8]
  PIN top_W6BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 268.600000 0.700000 268.980000 ;
    END
  END top_W6BEG[7]
  PIN top_W6BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.8844 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.712 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 267.380000 0.700000 267.760000 ;
    END
  END top_W6BEG[6]
  PIN top_W6BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 266.160000 0.700000 266.540000 ;
    END
  END top_W6BEG[5]
  PIN top_W6BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.1264 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.336 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 264.330000 0.700000 264.710000 ;
    END
  END top_W6BEG[4]
  PIN top_W6BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 263.110000 0.700000 263.490000 ;
    END
  END top_W6BEG[3]
  PIN top_W6BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.1604 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.184 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 261.280000 0.700000 261.660000 ;
    END
  END top_W6BEG[2]
  PIN top_W6BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 260.060000 0.700000 260.440000 ;
    END
  END top_W6BEG[1]
  PIN top_W6BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 258.230000 0.700000 258.610000 ;
    END
  END top_W6BEG[0]
  PIN top_W1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.228 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.016 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 15.2142 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 59.418 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.446055 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 60.6357 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 326.208 LAYER met4  ;
    ANTENNAGATEAREA 2.1837 LAYER met4  ;
    ANTENNAMAXAREACAR 73.3055 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 384.015 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.07799 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 209.430000 200.100000 209.810000 ;
    END
  END top_W1END[3]
  PIN top_W1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 13.1974 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 70.848 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 46.8374 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 226.879 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.394295 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 57.48 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 308.432 LAYER met4  ;
    ANTENNAGATEAREA 2.1837 LAYER met4  ;
    ANTENNAMAXAREACAR 73.1597 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 368.122 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.967925 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 207.600000 200.100000 207.980000 ;
    END
  END top_W1END[2]
  PIN top_W1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 13.1044 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 70.352 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 40.4555 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 194.313 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.446055 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 48.9879 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 263.616 LAYER met4  ;
    ANTENNAGATEAREA 1.8657 LAYER met4  ;
    ANTENNAMAXAREACAR 78.8472 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 408.851 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.47107 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 206.380000 200.100000 206.760000 ;
    END
  END top_W1END[1]
  PIN top_W1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 9.412 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 50.184 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 26.4035 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 120.929 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 70.3074 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 375.904 LAYER met4  ;
    ANTENNAGATEAREA 1.7067 LAYER met4  ;
    ANTENNAMAXAREACAR 74.5681 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 381.57 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 205.160000 200.100000 205.540000 ;
    END
  END top_W1END[0]
  PIN top_W2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 23.5842 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 126.248 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.8132 LAYER met3  ;
    ANTENNAMAXAREACAR 28.9915 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 144.261 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.354037 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 221.020000 200.100000 221.400000 ;
    END
  END top_W2MID[7]
  PIN top_W2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 24.0027 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 128.96 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6735 LAYER met3  ;
    ANTENNAMAXAREACAR 79.2324 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 402.779 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.382662 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 219.800000 200.100000 220.180000 ;
    END
  END top_W2MID[6]
  PIN top_W2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.67 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 169.36 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.5024 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 9.424 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8325 LAYER met4  ;
    ANTENNAMAXAREACAR 38.847 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 190.698 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.732075 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 217.970000 200.100000 218.350000 ;
    END
  END top_W2MID[5]
  PIN top_W2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 24.9742 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 134.128 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 9.975 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 55.552 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6735 LAYER met4  ;
    ANTENNAMAXAREACAR 69.6969 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 356.295 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.872265 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 216.750000 200.100000 217.130000 ;
    END
  END top_W2MID[4]
  PIN top_W2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 43.3126 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 230.992 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 22.9776 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 123.488 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8325 LAYER met4  ;
    ANTENNAMAXAREACAR 42.3712 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 223.049 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.07583 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 215.530000 200.100000 215.910000 ;
    END
  END top_W2MID[3]
  PIN top_W2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.6542 LAYER met3  ;
    ANTENNAMAXAREACAR 17.909 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 71.0377 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.347451 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 213.700000 200.100000 214.080000 ;
    END
  END top_W2MID[2]
  PIN top_W2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 26.2692 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 141.048 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8325 LAYER met3  ;
    ANTENNAMAXAREACAR 51.7533 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 264.223 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.512828 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 212.480000 200.100000 212.860000 ;
    END
  END top_W2MID[1]
  PIN top_W2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.2356 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 17.248 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 4.0806 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 22.704 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6735 LAYER met4  ;
    ANTENNAMAXAREACAR 28.7225 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 140.262 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.583562 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 210.650000 200.100000 211.030000 ;
    END
  END top_W2MID[0]
  PIN top_W2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 6.4593 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 34.44 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.6542 LAYER met3  ;
    ANTENNAMAXAREACAR 27.8972 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 126.422 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.508654 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 233.220000 200.100000 233.600000 ;
    END
  END top_W2END[7]
  PIN top_W2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 26.0074 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 139.168 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 76.1484 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 382.934 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.394295 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 3.9858 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 21.728 LAYER met4  ;
    ANTENNAGATEAREA 0.7527 LAYER met4  ;
    ANTENNAMAXAREACAR 81.4437 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 411.801 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.574843 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 231.390000 200.100000 231.770000 ;
    END
  END top_W2END[6]
  PIN top_W2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 39.5778 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 211.552 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7527 LAYER met3  ;
    ANTENNAMAXAREACAR 76.744 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 382.87 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.449057 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 230.170000 200.100000 230.550000 ;
    END
  END top_W2END[5]
  PIN top_W2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 54.9132 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 293.336 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3095 LAYER met3  ;
    ANTENNAMAXAREACAR 62.1033 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 319.558 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.574843 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 228.950000 200.100000 229.330000 ;
    END
  END top_W2END[4]
  PIN top_W2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 26.6901 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 143.288 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1505 LAYER met3  ;
    ANTENNAMAXAREACAR 64.911 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 325.817 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.548637 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 227.120000 200.100000 227.500000 ;
    END
  END top_W2END[3]
  PIN top_W2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 15.991 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 85.752 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9117 LAYER met3  ;
    ANTENNAMAXAREACAR 43.4562 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 204.215 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.454893 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.0338 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 5.984 LAYER met4  ;
    ANTENNAGATEAREA 1.3887 LAYER met4  ;
    ANTENNAMAXAREACAR 44.2006 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 208.524 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.632495 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 225.900000 200.100000 226.280000 ;
    END
  END top_W2END[2]
  PIN top_W2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 29.1784 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 156.08 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 73.9227 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 374.561 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.394295 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 4.7178 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 25.632 LAYER met4  ;
    ANTENNAGATEAREA 1.3887 LAYER met4  ;
    ANTENNAMAXAREACAR 77.32 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 393.018 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.758281 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 224.070000 200.100000 224.450000 ;
    END
  END top_W2END[1]
  PIN top_W2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 15.2904 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 82.024 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5145 LAYER met3  ;
    ANTENNAMAXAREACAR 64.6037 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 327.525 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.401016 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 222.850000 200.100000 223.230000 ;
    END
  END top_W2END[0]
  PIN top_WW4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.3166 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 33.68 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 3.705 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 22.112 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 31.3257 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 175.415 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 257.010000 200.100000 257.390000 ;
    END
  END top_WW4END[15]
  PIN top_WW4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9754 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 21.664 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.0514 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 12.352 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 43.4122 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 229.023 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 255.180000 200.100000 255.560000 ;
    END
  END top_WW4END[14]
  PIN top_WW4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 48.4486 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 258.384 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.2954 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.32 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 19.8463 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 109.562 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 253.960000 200.100000 254.340000 ;
    END
  END top_WW4END[13]
  PIN top_WW4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 29.353 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 157.016 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 9.4116 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 51.136 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 125.564 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 669.298 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 252.740000 200.100000 253.120000 ;
    END
  END top_WW4END[12]
  PIN top_WW4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 44.8204 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 239.504 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.2954 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.32 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 18.9969 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 105.038 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 250.910000 200.100000 251.290000 ;
    END
  END top_WW4END[11]
  PIN top_WW4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 46.1104 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 246.384 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.0676 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 11.968 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 21.9781 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 117.847 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 249.690000 200.100000 250.070000 ;
    END
  END top_WW4END[10]
  PIN top_WW4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 45.5344 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 243.312 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 17.7003 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 95.6947 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 247.860000 200.100000 248.240000 ;
    END
  END top_WW4END[9]
  PIN top_WW4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.849 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.328 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.5122 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 15.28 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 28.7415 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 159.98 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 246.640000 200.100000 247.020000 ;
    END
  END top_WW4END[8]
  PIN top_WW4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.1384 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 65.2 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 12.6174 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 68.704 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 75.1761 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 403.776 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 244.810000 200.100000 245.190000 ;
    END
  END top_WW4END[7]
  PIN top_WW4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 48.9334 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 261.44 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 3.1254 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 18.08 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 30.7415 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 168.621 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 243.590000 200.100000 243.970000 ;
    END
  END top_WW4END[6]
  PIN top_WW4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.3194 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 12.832 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 4.4916 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 27.248 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 104.758 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 553.288 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 242.370000 200.100000 242.750000 ;
    END
  END top_WW4END[5]
  PIN top_WW4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.8304 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 90.224 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 8.1384 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 44.816 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 67.2127 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 360.3 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 240.540000 200.100000 240.920000 ;
    END
  END top_WW4END[4]
  PIN top_WW4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 15.654 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 84.424 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9117 LAYER met3  ;
    ANTENNAMAXAREACAR 53.1895 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 267.061 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 239.320000 200.100000 239.700000 ;
    END
  END top_WW4END[3]
  PIN top_WW4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 45.4086 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 242.624 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 120.041 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 617.361 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.12 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.57833 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 18.1554 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 98.24 LAYER met4  ;
    ANTENNAGATEAREA 0.9117 LAYER met4  ;
    ANTENNAMAXAREACAR 139.954 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 725.116 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 237.490000 200.100000 237.870000 ;
    END
  END top_WW4END[2]
  PIN top_WW4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9936 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.624 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 4.6296 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 25.632 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9117 LAYER met4  ;
    ANTENNAMAXAREACAR 41.3405 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 206.341 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.501893 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 236.270000 200.100000 236.650000 ;
    END
  END top_WW4END[1]
  PIN top_WW4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 17.9134 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 96 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 66.5349 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 328.556 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.446055 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.1318 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 11.84 LAYER met4  ;
    ANTENNAGATEAREA 0.9117 LAYER met4  ;
    ANTENNAMAXAREACAR 68.8731 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 341.543 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.490985 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 234.440000 200.100000 234.820000 ;
    END
  END top_WW4END[0]
  PIN top_W6END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 20.038 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 107.336 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.1766 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 7.216 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 70.9018 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 368.239 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 274.700000 200.100000 275.080000 ;
    END
  END top_W6END[11]
  PIN top_W6END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 51.3466 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 273.84 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.3356 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.064 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 21.2758 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 115.394 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 273.480000 200.100000 273.860000 ;
    END
  END top_W6END[10]
  PIN top_W6END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 40.7416 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 217.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.3356 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.064 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 64.4804 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 346.392 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 271.650000 200.100000 272.030000 ;
    END
  END top_W6END[9]
  PIN top_W6END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 51.0274 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 272.608 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.9696 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 6.112 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 18.2331 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 98.2799 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 270.430000 200.100000 270.810000 ;
    END
  END top_W6END[8]
  PIN top_W6END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.468 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 168.296 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.3356 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.064 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 56.5186 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 304.168 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 268.600000 200.100000 268.980000 ;
    END
  END top_W6END[7]
  PIN top_W6END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5796 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.416 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.0514 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 12.352 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 37.943 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 204.122 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 267.380000 200.100000 267.760000 ;
    END
  END top_W6END[6]
  PIN top_W6END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.5216 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 45.44 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 3.8334 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 21.856 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 26.0224 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 143.802 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 266.160000 200.100000 266.540000 ;
    END
  END top_W6END[5]
  PIN top_W6END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.9166 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 68.88 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.631 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 16.384 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 23.2804 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 133.476 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 264.330000 200.100000 264.710000 ;
    END
  END top_W6END[4]
  PIN top_W6END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 43.954 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 234.888 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.3356 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.064 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 15.0779 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 83.598 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 263.110000 200.100000 263.490000 ;
    END
  END top_W6END[3]
  PIN top_W6END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 54.3076 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 289.632 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.2954 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.32 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 24.0631 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 132.249 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 261.280000 200.100000 261.660000 ;
    END
  END top_W6END[2]
  PIN top_W6END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 20.0494 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 107.392 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 60.3874 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 299.884 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.394295 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 12.1971 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 66.928 LAYER met4  ;
    ANTENNAGATEAREA 2.0247 LAYER met4  ;
    ANTENNAMAXAREACAR 66.4115 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 332.94 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 260.060000 200.100000 260.440000 ;
    END
  END top_W6END[1]
  PIN top_W6END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 22.822 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 122.184 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 65.0904 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 324.838 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.446055 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.6678 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.032 LAYER met4  ;
    ANTENNAGATEAREA 1.8657 LAYER met4  ;
    ANTENNAMAXAREACAR 65.4483 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 326.999 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.854368 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 258.230000 200.100000 258.610000 ;
    END
  END top_W6END[0]
  PIN bot_E1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.2504 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.664 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 80.720000 200.100000 81.100000 ;
    END
  END bot_E1BEG[3]
  PIN bot_E1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.9404 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.344 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 79.500000 200.100000 79.880000 ;
    END
  END bot_E1BEG[2]
  PIN bot_E1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 77.670000 200.100000 78.050000 ;
    END
  END bot_E1BEG[1]
  PIN bot_E1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 17.7084 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 94.44 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 76.450000 200.100000 76.830000 ;
    END
  END bot_E1BEG[0]
  PIN bot_E2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 92.920000 200.100000 93.300000 ;
    END
  END bot_E2BEG[7]
  PIN bot_E2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 91.700000 200.100000 92.080000 ;
    END
  END bot_E2BEG[6]
  PIN bot_E2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.6414 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.568 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 89.870000 200.100000 90.250000 ;
    END
  END bot_E2BEG[5]
  PIN bot_E2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 88.650000 200.100000 89.030000 ;
    END
  END bot_E2BEG[4]
  PIN bot_E2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 86.820000 200.100000 87.200000 ;
    END
  END bot_E2BEG[3]
  PIN bot_E2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.9884 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.6 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 85.600000 200.100000 85.980000 ;
    END
  END bot_E2BEG[2]
  PIN bot_E2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 83.770000 200.100000 84.150000 ;
    END
  END bot_E2BEG[1]
  PIN bot_E2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 82.550000 200.100000 82.930000 ;
    END
  END bot_E2BEG[0]
  PIN bot_E2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 105.120000 200.100000 105.500000 ;
    END
  END bot_E2BEGb[7]
  PIN bot_E2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 103.290000 200.100000 103.670000 ;
    END
  END bot_E2BEGb[6]
  PIN bot_E2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.6784 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 14.28 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 102.070000 200.100000 102.450000 ;
    END
  END bot_E2BEGb[5]
  PIN bot_E2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 100.240000 200.100000 100.620000 ;
    END
  END bot_E2BEGb[4]
  PIN bot_E2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.5744 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.392 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 99.020000 200.100000 99.400000 ;
    END
  END bot_E2BEGb[3]
  PIN bot_E2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 97.190000 200.100000 97.570000 ;
    END
  END bot_E2BEGb[2]
  PIN bot_E2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 95.970000 200.100000 96.350000 ;
    END
  END bot_E2BEGb[1]
  PIN bot_E2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 94.140000 200.100000 94.520000 ;
    END
  END bot_E2BEGb[0]
  PIN bot_EE4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.1264 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.336 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 128.910000 200.100000 129.290000 ;
    END
  END bot_EE4BEG[15]
  PIN bot_EE4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 127.080000 200.100000 127.460000 ;
    END
  END bot_EE4BEG[14]
  PIN bot_EE4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.6444 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 19.432 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 125.860000 200.100000 126.240000 ;
    END
  END bot_EE4BEG[13]
  PIN bot_EE4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 124.030000 200.100000 124.410000 ;
    END
  END bot_EE4BEG[12]
  PIN bot_EE4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.9884 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.6 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 122.810000 200.100000 123.190000 ;
    END
  END bot_EE4BEG[11]
  PIN bot_EE4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 121.590000 200.100000 121.970000 ;
    END
  END bot_EE4BEG[10]
  PIN bot_EE4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 119.760000 200.100000 120.140000 ;
    END
  END bot_EE4BEG[9]
  PIN bot_EE4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 118.540000 200.100000 118.920000 ;
    END
  END bot_EE4BEG[8]
  PIN bot_EE4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.1234 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.32 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 116.710000 200.100000 117.090000 ;
    END
  END bot_EE4BEG[7]
  PIN bot_EE4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.5744 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.392 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 115.490000 200.100000 115.870000 ;
    END
  END bot_EE4BEG[6]
  PIN bot_EE4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 113.660000 200.100000 114.040000 ;
    END
  END bot_EE4BEG[5]
  PIN bot_EE4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.8504 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.864 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 112.440000 200.100000 112.820000 ;
    END
  END bot_EE4BEG[4]
  PIN bot_EE4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 110.610000 200.100000 110.990000 ;
    END
  END bot_EE4BEG[3]
  PIN bot_EE4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 109.390000 200.100000 109.770000 ;
    END
  END bot_EE4BEG[2]
  PIN bot_EE4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.7124 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.128 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 107.560000 200.100000 107.940000 ;
    END
  END bot_EE4BEG[1]
  PIN bot_EE4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 106.340000 200.100000 106.720000 ;
    END
  END bot_EE4BEG[0]
  PIN bot_E6BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 146.600000 200.100000 146.980000 ;
    END
  END bot_E6BEG[11]
  PIN bot_E6BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.1604 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.184 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 145.380000 200.100000 145.760000 ;
    END
  END bot_E6BEG[10]
  PIN bot_E6BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 143.550000 200.100000 143.930000 ;
    END
  END bot_E6BEG[9]
  PIN bot_E6BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 142.330000 200.100000 142.710000 ;
    END
  END bot_E6BEG[8]
  PIN bot_E6BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 140.500000 200.100000 140.880000 ;
    END
  END bot_E6BEG[7]
  PIN bot_E6BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 139.280000 200.100000 139.660000 ;
    END
  END bot_E6BEG[6]
  PIN bot_E6BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.1604 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.184 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 137.450000 200.100000 137.830000 ;
    END
  END bot_E6BEG[5]
  PIN bot_E6BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.8504 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.864 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 136.230000 200.100000 136.610000 ;
    END
  END bot_E6BEG[4]
  PIN bot_E6BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.2504 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.664 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 135.010000 200.100000 135.390000 ;
    END
  END bot_E6BEG[3]
  PIN bot_E6BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 133.180000 200.100000 133.560000 ;
    END
  END bot_E6BEG[2]
  PIN bot_E6BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.2984 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.92 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 131.960000 200.100000 132.340000 ;
    END
  END bot_E6BEG[1]
  PIN bot_E6BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 130.130000 200.100000 130.510000 ;
    END
  END bot_E6BEG[0]
  PIN bot_E1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.6596 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 14.176 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 25.4658 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 138.64 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.1837 LAYER met4  ;
    ANTENNAMAXAREACAR 56.5199 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 303.243 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.07799 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 80.720000 0.700000 81.100000 ;
    END
  END bot_E1END[3]
  PIN bot_E1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 26.564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 142.128 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.0707 LAYER met3  ;
    ANTENNAMAXAREACAR 54.0387 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 269.415 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.472705 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 19.9614 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 107.872 LAYER met4  ;
    ANTENNAGATEAREA 2.1837 LAYER met4  ;
    ANTENNAMAXAREACAR 63.1798 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 318.814 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.07799 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 79.500000 0.700000 79.880000 ;
    END
  END bot_E1END[2]
  PIN bot_E1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 30.0145 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 161.48 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2297 LAYER met3  ;
    ANTENNAMAXAREACAR 41.6061 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 198.726 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.858943 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 28.8195 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 154.64 LAYER met4  ;
    ANTENNAGATEAREA 1.8657 LAYER met4  ;
    ANTENNAMAXAREACAR 57.0531 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 281.612 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.858943 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 77.670000 0.700000 78.050000 ;
    END
  END bot_E1END[1]
  PIN bot_E1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 9.0648 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 49.264 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7527 LAYER met3  ;
    ANTENNAMAXAREACAR 36.4654 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 179.34 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.769494 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.1558 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 11.968 LAYER met4  ;
    ANTENNAGATEAREA 1.8657 LAYER met4  ;
    ANTENNAMAXAREACAR 45.4106 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 225.994 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.769494 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 76.450000 0.700000 76.830000 ;
    END
  END bot_E1END[0]
  PIN bot_E2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 22.9264 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 122.736 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 15.807 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 86.656 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8325 LAYER met4  ;
    ANTENNAMAXAREACAR 49.9388 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 256.266 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.09371 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 92.920000 0.700000 93.300000 ;
    END
  END bot_E2MID[7]
  PIN bot_E2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.435 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.12 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 20.199 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 110.08 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8325 LAYER met4  ;
    ANTENNAMAXAREACAR 78.0234 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 408.76 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.47107 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 91.700000 0.700000 92.080000 ;
    END
  END bot_E2MID[6]
  PIN bot_E2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 25.1248 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 134.936 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.636 LAYER met3  ;
    ANTENNAMAXAREACAR 64.0445 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 325.996 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.51195 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 8.9478 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 50.544 LAYER met4  ;
    ANTENNAGATEAREA 0.8325 LAYER met4  ;
    ANTENNAMAXAREACAR 74.7926 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 386.71 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 89.870000 0.700000 90.250000 ;
    END
  END bot_E2MID[5]
  PIN bot_E2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.3809 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 77.52 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.477 LAYER met3  ;
    ANTENNAMAXAREACAR 67.8648 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 339.99 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.857862 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.6374 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 10.144 LAYER met4  ;
    ANTENNAGATEAREA 0.6735 LAYER met4  ;
    ANTENNAMAXAREACAR 70.296 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 355.051 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.857862 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 88.650000 0.700000 89.030000 ;
    END
  END bot_E2MID[4]
  PIN bot_E2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 32.6044 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 174.352 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.636 LAYER met3  ;
    ANTENNAMAXAREACAR 100.257 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 509.442 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.794969 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.5186 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 9.04 LAYER met4  ;
    ANTENNAGATEAREA 0.8325 LAYER met4  ;
    ANTENNAMAXAREACAR 102.081 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 520.301 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.794969 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 86.820000 0.700000 87.200000 ;
    END
  END bot_E2MID[3]
  PIN bot_E2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.3422 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 168.104 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6735 LAYER met3  ;
    ANTENNAMAXAREACAR 107.554 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 545.036 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.774004 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 85.600000 0.700000 85.980000 ;
    END
  END bot_E2MID[2]
  PIN bot_E2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 58.9011 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 315.08 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8325 LAYER met3  ;
    ANTENNAMAXAREACAR 88.114 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 457.753 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.574843 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 83.770000 0.700000 84.150000 ;
    END
  END bot_E2MID[1]
  PIN bot_E2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 26.1882 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 140.616 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8325 LAYER met3  ;
    ANTENNAMAXAREACAR 54.0247 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 271.651 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.590566 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 82.550000 0.700000 82.930000 ;
    END
  END bot_E2MID[0]
  PIN bot_E2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 9.2419 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 49.752 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5937 LAYER met3  ;
    ANTENNAMAXAREACAR 35.9043 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 167.253 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.354407 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.3052 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 14.176 LAYER met4  ;
    ANTENNAGATEAREA 1.2297 LAYER met4  ;
    ANTENNAMAXAREACAR 39.8034 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 201.366 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.695388 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 105.120000 0.700000 105.500000 ;
    END
  END bot_E2END[7]
  PIN bot_E2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 48.8626 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 261.048 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2297 LAYER met3  ;
    ANTENNAMAXAREACAR 52.2472 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 255.999 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.607371 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 6.3408 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 34.288 LAYER met4  ;
    ANTENNAGATEAREA 1.3887 LAYER met4  ;
    ANTENNAMAXAREACAR 56.8132 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 280.69 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 103.290000 0.700000 103.670000 ;
    END
  END bot_E2END[6]
  PIN bot_E2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.5226 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 24.112 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 22.6758 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 121.408 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3887 LAYER met4  ;
    ANTENNAMAXAREACAR 43.9969 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 223.114 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.870942 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 102.070000 0.700000 102.450000 ;
    END
  END bot_E2END[5]
  PIN bot_E2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 9.0536 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 48.744 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7527 LAYER met3  ;
    ANTENNAMAXAREACAR 46.7645 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 219.053 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.677348 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 3.5316 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 19.776 LAYER met4  ;
    ANTENNAGATEAREA 1.2297 LAYER met4  ;
    ANTENNAMAXAREACAR 49.6364 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 235.135 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 100.240000 0.700000 100.620000 ;
    END
  END bot_E2END[4]
  PIN bot_E2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 37.4332 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 200.096 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2297 LAYER met3  ;
    ANTENNAMAXAREACAR 68.1607 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 343.197 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.665023 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 8.1066 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 44.176 LAYER met4  ;
    ANTENNAGATEAREA 1.7067 LAYER met4  ;
    ANTENNAMAXAREACAR 72.9106 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 369.081 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 99.020000 0.700000 99.400000 ;
    END
  END bot_E2END[3]
  PIN bot_E2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 26.3764 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 141.136 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 71.2696 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 358.79 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.512537 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.6166 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 14.896 LAYER met4  ;
    ANTENNAGATEAREA 1.5477 LAYER met4  ;
    ANTENNAMAXAREACAR 72.9603 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 368.415 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.07799 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 97.190000 0.700000 97.570000 ;
    END
  END bot_E2END[2]
  PIN bot_E2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 7.7172 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 41.624 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.0707 LAYER met3  ;
    ANTENNAMAXAREACAR 22.0972 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 106.319 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.449057 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 95.970000 0.700000 96.350000 ;
    END
  END bot_E2END[1]
  PIN bot_E2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.366 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.752 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 16.1304 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 63.8567 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.394295 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 14.4888 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 77.744 LAYER met4  ;
    ANTENNAGATEAREA 1.0707 LAYER met4  ;
    ANTENNAMAXAREACAR 70.8943 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 359.58 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.590566 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 94.140000 0.700000 94.520000 ;
    END
  END bot_E2END[0]
  PIN bot_EE4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 44.6086 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 237.904 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.3356 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.064 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 28.7481 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 153.7 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 128.910000 0.700000 129.290000 ;
    END
  END bot_EE4END[15]
  PIN bot_EE4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 43.933 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 234.776 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.3356 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.064 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 33.972 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 175.7 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 127.080000 0.700000 127.460000 ;
    END
  END bot_EE4END[14]
  PIN bot_EE4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.4766 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 13.2 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 4.095 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 24.192 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 40.0768 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 221.069 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 125.860000 0.700000 126.240000 ;
    END
  END bot_EE4END[13]
  PIN bot_EE4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 39.7624 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 212.528 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.5186 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 9.04 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 26.4316 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 142.336 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 124.030000 0.700000 124.410000 ;
    END
  END bot_EE4END[12]
  PIN bot_EE4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 15.3496 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 81.856 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 7.3344 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 40.528 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 59.1537 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 312.748 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 122.810000 0.700000 123.190000 ;
    END
  END bot_EE4END[11]
  PIN bot_EE4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 51.982 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 277.704 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.3356 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.064 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 25.7084 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 133.186 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 121.590000 0.700000 121.970000 ;
    END
  END bot_EE4END[10]
  PIN bot_EE4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 55.3954 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 295.904 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.1526 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 7.088 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 19.5313 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 106.712 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 119.760000 0.700000 120.140000 ;
    END
  END bot_EE4END[9]
  PIN bot_EE4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 42.4906 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 226.608 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 24.0448 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 129.405 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 118.540000 0.700000 118.920000 ;
    END
  END bot_EE4END[8]
  PIN bot_EE4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 36.163 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 193.336 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.3052 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 14.176 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 29.345 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 163.216 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 116.710000 0.700000 117.090000 ;
    END
  END bot_EE4END[7]
  PIN bot_EE4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 34.8154 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 186.144 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.1462 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 13.328 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 38.8097 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 208.804 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 115.490000 0.700000 115.870000 ;
    END
  END bot_EE4END[6]
  PIN bot_EE4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 35.014 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 187.208 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.5186 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 9.04 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 20.4483 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 111.735 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 113.660000 0.700000 114.040000 ;
    END
  END bot_EE4END[5]
  PIN bot_EE4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.7896 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.536 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.4882 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 15.152 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 25.913 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 145.476 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 112.440000 0.700000 112.820000 ;
    END
  END bot_EE4END[4]
  PIN bot_EE4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7527 LAYER met3  ;
    ANTENNAMAXAREACAR 25.1956 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 106.992 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.376412 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 110.610000 0.700000 110.990000 ;
    END
  END bot_EE4END[3]
  PIN bot_EE4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 25.0384 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 134 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 75.404 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 378.091 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.446055 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.6678 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.032 LAYER met4  ;
    ANTENNAGATEAREA 0.9117 LAYER met4  ;
    ANTENNAMAXAREACAR 76.1364 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 382.513 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.774004 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 109.390000 0.700000 109.770000 ;
    END
  END bot_EE4END[2]
  PIN bot_EE4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.4096 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 34.176 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 6.9138 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 37.344 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9117 LAYER met4  ;
    ANTENNAMAXAREACAR 35.7858 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 176.531 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.411019 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 107.560000 0.700000 107.940000 ;
    END
  END bot_EE4END[1]
  PIN bot_EE4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 15.7311 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 84.36 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9117 LAYER met3  ;
    ANTENNAMAXAREACAR 46.8763 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 231.533 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.548637 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 106.340000 0.700000 106.720000 ;
    END
  END bot_EE4END[0]
  PIN bot_E6END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 52.2916 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 278.88 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.1526 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 7.088 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 23.1532 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 124.361 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 146.600000 0.700000 146.980000 ;
    END
  END bot_E6END[11]
  PIN bot_E6END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 52.2274 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 279.008 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.3356 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.064 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 25.6865 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 137.69 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 145.380000 0.700000 145.760000 ;
    END
  END bot_E6END[10]
  PIN bot_E6END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 17.578 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 94.216 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 4.6938 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 25.504 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 93.6555 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 497.425 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 143.550000 0.700000 143.930000 ;
    END
  END bot_E6END[9]
  PIN bot_E6END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 42.1246 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 224.656 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.2954 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.32 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 58.7888 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 317.384 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 142.330000 0.700000 142.710000 ;
    END
  END bot_E6END[8]
  PIN bot_E6END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 51.0496 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 272.256 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.9696 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 6.112 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 25.8316 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 133.064 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 140.500000 0.700000 140.880000 ;
    END
  END bot_E6END[7]
  PIN bot_E6END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 42.1246 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 224.656 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.2954 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.32 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 57.3135 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 308.438 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 139.280000 0.700000 139.660000 ;
    END
  END bot_E6END[6]
  PIN bot_E6END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.7014 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 41.536 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.8204 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 11.12 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 19.1186 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 106.025 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 137.450000 0.700000 137.830000 ;
    END
  END bot_E6END[5]
  PIN bot_E6END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 48.3346 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 257.776 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.3356 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.064 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 18.972 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 101.893 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 136.230000 0.700000 136.610000 ;
    END
  END bot_E6END[4]
  PIN bot_E6END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 47.479 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 253.688 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.3052 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 14.176 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 34.6672 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 184.763 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 135.010000 0.700000 135.390000 ;
    END
  END bot_E6END[3]
  PIN bot_E6END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 53.314 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 284.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.2954 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.32 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 15.5852 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 87.9033 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 133.180000 0.700000 133.560000 ;
    END
  END bot_E6END[2]
  PIN bot_E6END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 20.7795 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 112.696 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.3427 LAYER met3  ;
    ANTENNAMAXAREACAR 46.0527 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 224.148 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.590566 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 131.960000 0.700000 132.340000 ;
    END
  END bot_E6END[1]
  PIN bot_E6END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 17.5561 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 94.56 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.5477 LAYER met3  ;
    ANTENNAMAXAREACAR 43.5656 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 212.966 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.600688 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.4848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 3.056 LAYER met4  ;
    ANTENNAGATEAREA 2.3427 LAYER met4  ;
    ANTENNAMAXAREACAR 47.2482 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 239.428 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.625157 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 130.130000 0.700000 130.510000 ;
    END
  END bot_E6END[0]
  PIN bot_W1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.9204 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 20.904 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 9.350000 0.700000 9.730000 ;
    END
  END bot_W1BEG[3]
  PIN bot_W1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 7.520000 0.700000 7.900000 ;
    END
  END bot_W1BEG[2]
  PIN bot_W1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.9884 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.6 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 6.300000 0.700000 6.680000 ;
    END
  END bot_W1BEG[1]
  PIN bot_W1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 5.080000 0.700000 5.460000 ;
    END
  END bot_W1BEG[0]
  PIN bot_W2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 20.940000 0.700000 21.320000 ;
    END
  END bot_W2BEG[7]
  PIN bot_W2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 19.720000 0.700000 20.100000 ;
    END
  END bot_W2BEG[6]
  PIN bot_W2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 18.500000 0.700000 18.880000 ;
    END
  END bot_W2BEG[5]
  PIN bot_W2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.4024 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 12.808 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 16.670000 0.700000 17.050000 ;
    END
  END bot_W2BEG[4]
  PIN bot_W2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 15.450000 0.700000 15.830000 ;
    END
  END bot_W2BEG[3]
  PIN bot_W2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.2964 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.576 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 13.620000 0.700000 14.000000 ;
    END
  END bot_W2BEG[2]
  PIN bot_W2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 12.400000 0.700000 12.780000 ;
    END
  END bot_W2BEG[1]
  PIN bot_W2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 10.570000 0.700000 10.950000 ;
    END
  END bot_W2BEG[0]
  PIN bot_W2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 33.140000 0.700000 33.520000 ;
    END
  END bot_W2BEGb[7]
  PIN bot_W2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 31.920000 0.700000 32.300000 ;
    END
  END bot_W2BEGb[6]
  PIN bot_W2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 18.0414 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 96.216 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 30.090000 0.700000 30.470000 ;
    END
  END bot_W2BEGb[5]
  PIN bot_W2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 28.870000 0.700000 29.250000 ;
    END
  END bot_W2BEGb[4]
  PIN bot_W2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 27.040000 0.700000 27.420000 ;
    END
  END bot_W2BEGb[3]
  PIN bot_W2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 18.5454 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 98.904 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 25.820000 0.700000 26.200000 ;
    END
  END bot_W2BEGb[2]
  PIN bot_W2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 23.990000 0.700000 24.370000 ;
    END
  END bot_W2BEGb[1]
  PIN bot_W2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 13.0704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 69.704 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 22.770000 0.700000 23.150000 ;
    END
  END bot_W2BEGb[0]
  PIN bot_WW4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.9504 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.064 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 56.930000 0.700000 57.310000 ;
    END
  END bot_WW4BEG[15]
  PIN bot_WW4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.1604 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.184 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 55.710000 0.700000 56.090000 ;
    END
  END bot_WW4BEG[14]
  PIN bot_WW4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 53.880000 0.700000 54.260000 ;
    END
  END bot_WW4BEG[13]
  PIN bot_WW4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.6104 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 24.584 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 52.660000 0.700000 53.040000 ;
    END
  END bot_WW4BEG[12]
  PIN bot_WW4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 50.830000 0.700000 51.210000 ;
    END
  END bot_WW4BEG[11]
  PIN bot_WW4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.8504 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.864 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 49.610000 0.700000 49.990000 ;
    END
  END bot_WW4BEG[10]
  PIN bot_WW4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 48.390000 0.700000 48.770000 ;
    END
  END bot_WW4BEG[9]
  PIN bot_WW4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.5744 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.392 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 46.560000 0.700000 46.940000 ;
    END
  END bot_WW4BEG[8]
  PIN bot_WW4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 45.340000 0.700000 45.720000 ;
    END
  END bot_WW4BEG[7]
  PIN bot_WW4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 43.510000 0.700000 43.890000 ;
    END
  END bot_WW4BEG[6]
  PIN bot_WW4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.8504 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.864 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 42.290000 0.700000 42.670000 ;
    END
  END bot_WW4BEG[5]
  PIN bot_WW4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 40.460000 0.700000 40.840000 ;
    END
  END bot_WW4BEG[4]
  PIN bot_WW4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.8844 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.712 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 39.240000 0.700000 39.620000 ;
    END
  END bot_WW4BEG[3]
  PIN bot_WW4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 37.410000 0.700000 37.790000 ;
    END
  END bot_WW4BEG[2]
  PIN bot_WW4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.0224 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.448 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 36.190000 0.700000 36.570000 ;
    END
  END bot_WW4BEG[1]
  PIN bot_WW4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 34.360000 0.700000 34.740000 ;
    END
  END bot_WW4BEG[0]
  PIN bot_W6BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.6554 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 24.824 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 75.230000 0.700000 75.610000 ;
    END
  END bot_W6BEG[11]
  PIN bot_W6BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 73.400000 0.700000 73.780000 ;
    END
  END bot_W6BEG[10]
  PIN bot_W6BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.0224 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.448 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 72.180000 0.700000 72.560000 ;
    END
  END bot_W6BEG[9]
  PIN bot_W6BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 70.350000 0.700000 70.730000 ;
    END
  END bot_W6BEG[8]
  PIN bot_W6BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 69.130000 0.700000 69.510000 ;
    END
  END bot_W6BEG[7]
  PIN bot_W6BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 67.300000 0.700000 67.680000 ;
    END
  END bot_W6BEG[6]
  PIN bot_W6BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.7124 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.128 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 66.080000 0.700000 66.460000 ;
    END
  END bot_W6BEG[5]
  PIN bot_W6BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 64.250000 0.700000 64.630000 ;
    END
  END bot_W6BEG[4]
  PIN bot_W6BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 63.030000 0.700000 63.410000 ;
    END
  END bot_W6BEG[3]
  PIN bot_W6BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 61.810000 0.700000 62.190000 ;
    END
  END bot_W6BEG[2]
  PIN bot_W6BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 59.980000 0.700000 60.360000 ;
    END
  END bot_W6BEG[1]
  PIN bot_W6BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 58.760000 0.700000 59.140000 ;
    END
  END bot_W6BEG[0]
  PIN bot_W1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 15.5194 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 83.232 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 70.7511 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 347.872 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.512537 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 19.9473 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 107.792 LAYER met4  ;
    ANTENNAGATEAREA 2.1837 LAYER met4  ;
    ANTENNAMAXAREACAR 79.8857 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 397.234 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 9.350000 200.100000 9.730000 ;
    END
  END bot_W1END[3]
  PIN bot_W1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 26.8662 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 143.752 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.1837 LAYER met3  ;
    ANTENNAMAXAREACAR 55.5789 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 275.147 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.656604 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 7.520000 200.100000 7.900000 ;
    END
  END bot_W1END[2]
  PIN bot_W1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 10.9252 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 59.2 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5937 LAYER met3  ;
    ANTENNAMAXAREACAR 58.5496 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 281.543 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 1.0353 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 15.1296 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 83.984 LAYER met4  ;
    ANTENNAGATEAREA 1.8657 LAYER met4  ;
    ANTENNAMAXAREACAR 66.6589 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 342.933 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.47107 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 6.300000 200.100000 6.680000 ;
    END
  END bot_W1END[1]
  PIN bot_W1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 7.2973 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 39.376 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5937 LAYER met3  ;
    ANTENNAMAXAREACAR 37.986 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 175.849 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.642217 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 14.4072 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 78.72 LAYER met4  ;
    ANTENNAGATEAREA 1.7067 LAYER met4  ;
    ANTENNAMAXAREACAR 73.7132 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 383.501 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 5.080000 200.100000 5.460000 ;
    END
  END bot_W1END[0]
  PIN bot_W2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1824 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.248 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 50.8229 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 254.893 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.872265 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 43.0128 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 229.872 LAYER met4  ;
    ANTENNAGATEAREA 0.8325 LAYER met4  ;
    ANTENNAMAXAREACAR 102.49 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 531.016 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.872265 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 20.940000 200.100000 21.320000 ;
    END
  END bot_W2MID[7]
  PIN bot_W2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3726 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.312 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 39.5568 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 213.792 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6735 LAYER met4  ;
    ANTENNAMAXAREACAR 78.8895 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 413.316 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 19.720000 200.100000 20.100000 ;
    END
  END bot_W2MID[6]
  PIN bot_W2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 38.3926 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 204.752 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 26.6475 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 143.056 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8325 LAYER met4  ;
    ANTENNAMAXAREACAR 54.081 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 276.418 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 18.500000 200.100000 18.880000 ;
    END
  END bot_W2MID[5]
  PIN bot_W2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5796 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.416 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 29.262 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 158.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6735 LAYER met4  ;
    ANTENNAMAXAREACAR 57.4538 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 305.483 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 16.670000 200.100000 17.050000 ;
    END
  END bot_W2MID[4]
  PIN bot_W2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7626 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.392 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 3.1896 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 17.952 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8325 LAYER met4  ;
    ANTENNAMAXAREACAR 30.9864 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 154.338 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.419367 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 15.450000 200.100000 15.830000 ;
    END
  END bot_W2MID[3]
  PIN bot_W2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 32.697 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 174.56 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 25.164 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 136.56 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6735 LAYER met4  ;
    ANTENNAMAXAREACAR 57.4799 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 298.164 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 13.620000 200.100000 14.000000 ;
    END
  END bot_W2MID[2]
  PIN bot_W2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 56.4972 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 302.264 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8325 LAYER met3  ;
    ANTENNAMAXAREACAR 88.8397 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 463.449 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.531572 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 12.400000 200.100000 12.780000 ;
    END
  END bot_W2MID[1]
  PIN bot_W2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5754 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.544 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8325 LAYER met3  ;
    ANTENNAMAXAREACAR 26.4422 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 125.957 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.512828 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 10.570000 200.100000 10.950000 ;
    END
  END bot_W2MID[0]
  PIN bot_W2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.1354 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 65.184 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 6.0132 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 33.952 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6735 LAYER met4  ;
    ANTENNAMAXAREACAR 78.1268 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 400.161 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.80021 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 33.140000 200.100000 33.520000 ;
    END
  END bot_W2END[7]
  PIN bot_W2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7527 LAYER met3  ;
    ANTENNAMAXAREACAR 18.394 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 73.1998 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.376412 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 31.920000 200.100000 32.300000 ;
    END
  END bot_W2END[6]
  PIN bot_W2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 21.4804 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 115.024 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 65.9972 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 328.624 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.446055 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 43.5696 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 233.312 LAYER met4  ;
    ANTENNAGATEAREA 0.7527 LAYER met4  ;
    ANTENNAMAXAREACAR 123.882 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 638.591 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.574843 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 30.090000 200.100000 30.470000 ;
    END
  END bot_W2END[5]
  PIN bot_W2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 42.7914 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 228.696 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3095 LAYER met3  ;
    ANTENNAMAXAREACAR 65.9604 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 333.568 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.495326 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 28.870000 200.100000 29.250000 ;
    END
  END bot_W2END[4]
  PIN bot_W2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 27.0652 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 145.28 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.795 LAYER met3  ;
    ANTENNAMAXAREACAR 68.3799 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 347.53 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.615723 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.5362 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 15.408 LAYER met4  ;
    ANTENNAGATEAREA 1.1505 LAYER met4  ;
    ANTENNAMAXAREACAR 70.5844 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 360.922 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.07799 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 27.040000 200.100000 27.420000 ;
    END
  END bot_W2END[3]
  PIN bot_W2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3887 LAYER met3  ;
    ANTENNAMAXAREACAR 27.9187 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 131.681 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.635093 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 25.820000 200.100000 26.200000 ;
    END
  END bot_W2END[2]
  PIN bot_W2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 37.899 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 203.064 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3887 LAYER met3  ;
    ANTENNAMAXAREACAR 46.5302 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 235.333 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.506709 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 23.990000 200.100000 24.370000 ;
    END
  END bot_W2END[1]
  PIN bot_W2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 37.5496 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 200.256 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6678 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.032 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5145 LAYER met4  ;
    ANTENNAMAXAREACAR 21.1082 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 100.756 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.620271 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 22.770000 200.100000 23.150000 ;
    END
  END bot_W2END[0]
  PIN bot_WW4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 43.225 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 231 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 13.2193 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 72.7684 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 56.930000 200.100000 57.310000 ;
    END
  END bot_WW4END[15]
  PIN bot_WW4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 52.9456 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 282.368 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 12.2372 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 66.3562 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 55.710000 200.100000 56.090000 ;
    END
  END bot_WW4END[14]
  PIN bot_WW4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 51.1414 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 273.216 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.9696 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 6.112 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 14.3308 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 78.8855 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 53.880000 200.100000 54.260000 ;
    END
  END bot_WW4END[13]
  PIN bot_WW4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 46.0606 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 245.648 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.3356 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.064 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 44.3069 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 238.392 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 52.660000 200.100000 53.040000 ;
    END
  END bot_WW4END[12]
  PIN bot_WW4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.3677 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 24.24 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 56.888 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 292.01 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.46514 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 50.830000 200.100000 51.210000 ;
    END
  END bot_WW4END[11]
  PIN bot_WW4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 37.0492 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 198.528 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.3258 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 2.208 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 30.2468 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 160.316 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 49.610000 200.100000 49.990000 ;
    END
  END bot_WW4END[10]
  PIN bot_WW4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.6016 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 19.2 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 3.1494 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 18.208 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 23.7237 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 131.41 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 48.390000 200.100000 48.770000 ;
    END
  END bot_WW4END[9]
  PIN bot_WW4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 48.9574 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 261.568 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.3356 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.064 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 22.8585 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 120.774 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 46.560000 200.100000 46.940000 ;
    END
  END bot_WW4END[8]
  PIN bot_WW4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 42.046 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 224.712 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.2954 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.32 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 23.9247 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 130.153 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 45.340000 200.100000 45.720000 ;
    END
  END bot_WW4END[7]
  PIN bot_WW4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 48.0736 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 256.384 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.6614 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 10.272 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 47.7104 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 258.041 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 43.510000 200.100000 43.890000 ;
    END
  END bot_WW4END[6]
  PIN bot_WW4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.4964 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 61.776 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 7.6698 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 41.376 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 49.9628 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 266.636 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 42.290000 200.100000 42.670000 ;
    END
  END bot_WW4END[5]
  PIN bot_WW4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1089 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.056 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 48.9267 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 242.636 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.46514 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 40.460000 200.100000 40.840000 ;
    END
  END bot_WW4END[4]
  PIN bot_WW4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.2863 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 28.632 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5937 LAYER met3  ;
    ANTENNAMAXAREACAR 22.0289 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 94.9344 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.642217 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 8.9508 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 48.208 LAYER met4  ;
    ANTENNAGATEAREA 0.9117 LAYER met4  ;
    ANTENNAMAXAREACAR 65.0182 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 332.668 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.716352 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 39.240000 200.100000 39.620000 ;
    END
  END bot_WW4END[3]
  PIN bot_WW4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 17.3392 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 93.408 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7527 LAYER met3  ;
    ANTENNAMAXAREACAR 52.2744 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 263.203 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.627985 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 5.9652 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 33.696 LAYER met4  ;
    ANTENNAGATEAREA 0.9117 LAYER met4  ;
    ANTENNAMAXAREACAR 58.8173 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 300.162 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 37.410000 200.100000 37.790000 ;
    END
  END bot_WW4END[2]
  PIN bot_WW4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 15.1743 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 81.368 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5937 LAYER met3  ;
    ANTENNAMAXAREACAR 38.6226 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 183.454 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.642217 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 17.6544 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 95.568 LAYER met4  ;
    ANTENNAGATEAREA 0.9117 LAYER met4  ;
    ANTENNAMAXAREACAR 57.9869 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 288.278 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 36.190000 200.100000 36.570000 ;
    END
  END bot_WW4END[1]
  PIN bot_WW4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 16.9968 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 91.12 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9117 LAYER met3  ;
    ANTENNAMAXAREACAR 61.754 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 309.93 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.42052 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 34.360000 200.100000 34.740000 ;
    END
  END bot_WW4END[0]
  PIN bot_W6END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 53.2804 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 284.624 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.9696 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 6.112 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 12.3949 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 68.5038 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 75.230000 200.100000 75.610000 ;
    END
  END bot_W6END[11]
  PIN bot_W6END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 41.29 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 220.68 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.4848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 3.056 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 29.1961 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 145.69 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 73.400000 200.100000 73.780000 ;
    END
  END bot_W6END[10]
  PIN bot_W6END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 53.8936 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 287.424 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.3356 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.064 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 18.7837 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 102.005 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 72.180000 200.100000 72.560000 ;
    END
  END bot_W6END[9]
  PIN bot_W6END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 26.2774 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 140.608 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 4.461 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 26.144 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 48.2417 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 265.242 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 70.350000 200.100000 70.730000 ;
    END
  END bot_W6END[8]
  PIN bot_W6END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.0104 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 27.184 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.265 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 14.432 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 48.9903 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 263.394 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 69.130000 200.100000 69.510000 ;
    END
  END bot_W6END[7]
  PIN bot_W6END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.975 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 171 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.9696 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 6.112 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 63.7069 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 334.728 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 67.300000 200.100000 67.680000 ;
    END
  END bot_W6END[6]
  PIN bot_W6END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.6424 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 35.888 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.9568 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 18.592 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 31.655 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 180.331 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 66.080000 200.100000 66.460000 ;
    END
  END bot_W6END[5]
  PIN bot_W6END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.7364 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 47.056 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.6212 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 10.528 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 27.512 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 152.784 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 64.250000 200.100000 64.630000 ;
    END
  END bot_W6END[4]
  PIN bot_W6END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 50.8444 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 271.632 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 3.4914 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 20.032 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 26.9567 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 147.399 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 63.030000 200.100000 63.410000 ;
    END
  END bot_W6END[3]
  PIN bot_W6END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.589 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 67.608 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.6614 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 10.272 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 29.0641 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 151.679 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 61.810000 200.100000 62.190000 ;
    END
  END bot_W6END[2]
  PIN bot_W6END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 33.2641 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 178.336 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.0707 LAYER met3  ;
    ANTENNAMAXAREACAR 54.2128 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 275.156 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.811363 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 3.0468 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 16.72 LAYER met4  ;
    ANTENNAGATEAREA 2.0247 LAYER met4  ;
    ANTENNAMAXAREACAR 55.7177 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 283.414 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.811363 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 59.980000 200.100000 60.360000 ;
    END
  END bot_W6END[1]
  PIN bot_W6END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.0884 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.6 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7527 LAYER met3  ;
    ANTENNAMAXAREACAR 26.9974 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 130.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.624206 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 13.5807 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 75.248 LAYER met4  ;
    ANTENNAGATEAREA 1.8657 LAYER met4  ;
    ANTENNAMAXAREACAR 34.2765 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 170.652 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 58.760000 200.100000 59.140000 ;
    END
  END bot_W6END[0]
  PIN bot_S1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.003 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.907 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 88.820000 0.000000 89.200000 0.700000 ;
    END
  END bot_S1BEG[3]
  PIN bot_S1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.3458 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.503 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 87.440000 0.000000 87.820000 0.700000 ;
    END
  END bot_S1BEG[2]
  PIN bot_S1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 7.3226 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 36.505 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 86.060000 0.000000 86.440000 0.700000 ;
    END
  END bot_S1BEG[1]
  PIN bot_S1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.965 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.599 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 84.220000 0.000000 84.600000 0.700000 ;
    END
  END bot_S1BEG[0]
  PIN bot_S2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.6386 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.085 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 113.200000 0.000000 113.580000 0.700000 ;
    END
  END bot_S2BEG[7]
  PIN bot_S2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.129 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.537 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 111.820000 0.000000 112.200000 0.700000 ;
    END
  END bot_S2BEG[6]
  PIN bot_S2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.2718 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.251 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 110.440000 0.000000 110.820000 0.700000 ;
    END
  END bot_S2BEG[5]
  PIN bot_S2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.8434 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.109 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 108.600000 0.000000 108.980000 0.700000 ;
    END
  END bot_S2BEG[4]
  PIN bot_S2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.9382 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.583 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 107.220000 0.000000 107.600000 0.700000 ;
    END
  END bot_S2BEG[3]
  PIN bot_S2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7338 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.561 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 105.840000 0.000000 106.220000 0.700000 ;
    END
  END bot_S2BEG[2]
  PIN bot_S2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.8434 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.109 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 104.000000 0.000000 104.380000 0.700000 ;
    END
  END bot_S2BEG[1]
  PIN bot_S2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.1766 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.775 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 102.620000 0.000000 103.000000 0.700000 ;
    END
  END bot_S2BEG[0]
  PIN bot_S2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.2886 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.335 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 101.240000 0.000000 101.620000 0.700000 ;
    END
  END bot_S2BEGb[7]
  PIN bot_S2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.8434 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.109 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 99.400000 0.000000 99.780000 0.700000 ;
    END
  END bot_S2BEGb[6]
  PIN bot_S2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.5742 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.763 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 98.020000 0.000000 98.400000 0.700000 ;
    END
  END bot_S2BEGb[5]
  PIN bot_S2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.2284 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.034 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 96.640000 0.000000 97.020000 0.700000 ;
    END
  END bot_S2BEGb[4]
  PIN bot_S2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.965 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.599 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 95.260000 0.000000 95.640000 0.700000 ;
    END
  END bot_S2BEGb[3]
  PIN bot_S2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7175 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.4265 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.2509 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 8.3538 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 45.024 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 93.420000 0.000000 93.800000 0.700000 ;
    END
  END bot_S2BEGb[2]
  PIN bot_S2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.6314 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.931 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 92.040000 0.000000 92.420000 0.700000 ;
    END
  END bot_S2BEGb[1]
  PIN bot_S2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.2928 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.356 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 90.660000 0.000000 91.040000 0.700000 ;
    END
  END bot_S2BEGb[0]
  PIN bot_S4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.9238 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.511 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 138.040000 0.000000 138.420000 0.700000 ;
    END
  END bot_S4BEG[15]
  PIN bot_S4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.6694 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.239 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 136.200000 0.000000 136.580000 0.700000 ;
    END
  END bot_S4BEG[14]
  PIN bot_S4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.2242 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.013 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 134.820000 0.000000 135.200000 0.700000 ;
    END
  END bot_S4BEG[13]
  PIN bot_S4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.1622 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.703 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 133.440000 0.000000 133.820000 0.700000 ;
    END
  END bot_S4BEG[12]
  PIN bot_S4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.2718 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.251 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 131.600000 0.000000 131.980000 0.700000 ;
    END
  END bot_S4BEG[11]
  PIN bot_S4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.8434 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.109 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 130.220000 0.000000 130.600000 0.700000 ;
    END
  END bot_S4BEG[10]
  PIN bot_S4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6321 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.9995 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.7518 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 20.48 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 128.840000 0.000000 129.220000 0.700000 ;
    END
  END bot_S4BEG[9]
  PIN bot_S4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.8434 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.109 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 127.000000 0.000000 127.380000 0.700000 ;
    END
  END bot_S4BEG[8]
  PIN bot_S4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.6862 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.323 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 125.620000 0.000000 126.000000 0.700000 ;
    END
  END bot_S4BEG[7]
  PIN bot_S4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.9862 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.823 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 124.240000 0.000000 124.620000 0.700000 ;
    END
  END bot_S4BEG[6]
  PIN bot_S4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.3362 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.573 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 122.400000 0.000000 122.780000 0.700000 ;
    END
  END bot_S4BEG[5]
  PIN bot_S4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.8434 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.109 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 121.020000 0.000000 121.400000 0.700000 ;
    END
  END bot_S4BEG[4]
  PIN bot_S4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.5574 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.679 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 119.640000 0.000000 120.020000 0.700000 ;
    END
  END bot_S4BEG[3]
  PIN bot_S4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.2242 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.013 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 117.800000 0.000000 118.180000 0.700000 ;
    END
  END bot_S4BEG[2]
  PIN bot_S4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7338 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.561 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 116.420000 0.000000 116.800000 0.700000 ;
    END
  END bot_S4BEG[1]
  PIN bot_S4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.8434 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.109 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 115.040000 0.000000 115.420000 0.700000 ;
    END
  END bot_S4BEG[0]
  PIN bot_SS4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6321 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.9995 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.2509 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 13.5018 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 72.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 162.420000 0.000000 162.800000 0.700000 ;
    END
  END bot_SS4BEG[15]
  PIN bot_SS4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.4482 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.133 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 160.580000 0.000000 160.960000 0.700000 ;
    END
  END bot_SS4BEG[14]
  PIN bot_SS4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.965 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.599 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 159.200000 0.000000 159.580000 0.700000 ;
    END
  END bot_SS4BEG[13]
  PIN bot_SS4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.2886 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.335 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 157.820000 0.000000 158.200000 0.700000 ;
    END
  END bot_SS4BEG[12]
  PIN bot_SS4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7814 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.799 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 155.980000 0.000000 156.360000 0.700000 ;
    END
  END bot_SS4BEG[11]
  PIN bot_SS4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.9382 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.583 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 154.600000 0.000000 154.980000 0.700000 ;
    END
  END bot_SS4BEG[10]
  PIN bot_SS4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.912 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.452 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 153.220000 0.000000 153.600000 0.700000 ;
    END
  END bot_SS4BEG[9]
  PIN bot_SS4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.965 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.599 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 151.380000 0.000000 151.760000 0.700000 ;
    END
  END bot_SS4BEG[8]
  PIN bot_SS4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6965 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.3215 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.4758 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 19.008 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 150.000000 0.000000 150.380000 0.700000 ;
    END
  END bot_SS4BEG[7]
  PIN bot_SS4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.5098 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.441 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 148.620000 0.000000 149.000000 0.700000 ;
    END
  END bot_SS4BEG[6]
  PIN bot_SS4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.2578 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.181 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 146.780000 0.000000 147.160000 0.700000 ;
    END
  END bot_SS4BEG[5]
  PIN bot_SS4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.465 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.217 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 145.400000 0.000000 145.780000 0.700000 ;
    END
  END bot_SS4BEG[4]
  PIN bot_SS4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.9722 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.753 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 144.020000 0.000000 144.400000 0.700000 ;
    END
  END bot_SS4BEG[3]
  PIN bot_SS4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.9914 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.849 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 142.640000 0.000000 143.020000 0.700000 ;
    END
  END bot_SS4BEG[2]
  PIN bot_SS4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.3537 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.6605 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 140.800000 0.000000 141.180000 0.700000 ;
    END
  END bot_SS4BEG[1]
  PIN bot_SS4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7646 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.715 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 139.420000 0.000000 139.800000 0.700000 ;
    END
  END bot_SS4BEG[0]
  PIN bot_N1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.5223 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 27.4505 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 7.4404 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 40.144 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5937 LAYER met3  ;
    ANTENNAMAXAREACAR 22.3285 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 98.1479 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.458019 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 38.9565 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 208.704 LAYER met4  ;
    ANTENNAGATEAREA 2.0247 LAYER met4  ;
    ANTENNAMAXAREACAR 84.9495 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 428.084 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 9.240000 0.000000 9.620000 0.700000 ;
    END
  END bot_N1END[3]
  PIN bot_N1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.5009 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 31.8815 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7527 LAYER met2  ;
    ANTENNAMAXAREACAR 23.5135 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 107.771 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.517922 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.745 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.44 LAYER met3  ;
    ANTENNAGATEAREA 0.7527 LAYER met3  ;
    ANTENNAMAXAREACAR 24.5033 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 113.67 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.571064 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 15.5388 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 83.344 LAYER met4  ;
    ANTENNAGATEAREA 2.0247 LAYER met4  ;
    ANTENNAMAXAREACAR 58.8602 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 299.515 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.571064 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 7.860000 0.000000 8.240000 0.700000 ;
    END
  END bot_N1END[2]
  PIN bot_N1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.8816 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 23.968 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 21.6805 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 89.2604 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.354037 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 33.1026 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 177.936 LAYER met3  ;
    ANTENNAGATEAREA 1.0707 LAYER met3  ;
    ANTENNAMAXAREACAR 68.7327 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 345.803 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 1.00528 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 44.7756 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 239.264 LAYER met4  ;
    ANTENNAGATEAREA 2.0247 LAYER met4  ;
    ANTENNAMAXAREACAR 90.8474 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 463.976 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.00528 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 6.480000 0.000000 6.860000 0.700000 ;
    END
  END bot_N1END[1]
  PIN bot_N1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.7613 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.5275 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 13.0943 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 46.7 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.26202 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.161 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 27.992 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 24.9669 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 111.094 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.354037 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 32.7345 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 175.52 LAYER met4  ;
    ANTENNAGATEAREA 2.0247 LAYER met4  ;
    ANTENNAMAXAREACAR 76.5912 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 393.677 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.967925 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 5.100000 0.000000 5.480000 0.700000 ;
    END
  END bot_N1END[0]
  PIN bot_N2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2089 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.8835 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 92.4627 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 495.952 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.0247 LAYER met4  ;
    ANTENNAMAXAREACAR 114.307 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 592.5 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.32956 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 21.660000 0.000000 22.040000 0.700000 ;
    END
  END bot_N2MID[7]
  PIN bot_N2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1025 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.3515 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.09 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 73.8498 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 396.688 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.8657 LAYER met4  ;
    ANTENNAMAXAREACAR 96.2618 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 491.243 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.32956 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 20.280000 0.000000 20.660000 0.700000 ;
    END
  END bot_N2MID[6]
  PIN bot_N2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.1955 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.8165 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.3 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 39.4 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 67.3731 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 360.72 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.8657 LAYER met4  ;
    ANTENNAMAXAREACAR 80.4224 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 407.698 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 18.440000 0.000000 18.820000 0.700000 ;
    END
  END bot_N2MID[5]
  PIN bot_N2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.8711 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.1945 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.332 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 12.904 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 82.2408 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 440.96 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.8657 LAYER met4  ;
    ANTENNAMAXAREACAR 73.4307 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 376.457 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.632495 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 17.060000 0.000000 17.440000 0.700000 ;
    END
  END bot_N2MID[4]
  PIN bot_N2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8883 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.2805 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.883 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.176 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 91.005 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 487.712 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.0247 LAYER met4  ;
    ANTENNAMAXAREACAR 90.4535 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 465.691 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.02558 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 15.680000 0.000000 16.060000 0.700000 ;
    END
  END bot_N2MID[3]
  PIN bot_N2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1255 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.4565 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 16.774 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 89.928 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 30.2976 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 162.528 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.7067 LAYER met4  ;
    ANTENNAMAXAREACAR 74.4457 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 366.253 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.648174 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 13.840000 0.000000 14.220000 0.700000 ;
    END
  END bot_N2MID[2]
  PIN bot_N2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7175 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.4265 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.26895 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.832 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 84.2262 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 451.088 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.8657 LAYER met4  ;
    ANTENNAMAXAREACAR 83.3056 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 424.838 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.80021 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 12.460000 0.000000 12.840000 0.700000 ;
    END
  END bot_N2MID[1]
  PIN bot_N2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.6817 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.2475 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 16.4677 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 88.768 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2297 LAYER met3  ;
    ANTENNAMAXAREACAR 65.2299 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 322.039 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.562365 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 31.7856 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 170.464 LAYER met4  ;
    ANTENNAGATEAREA 2.0247 LAYER met4  ;
    ANTENNAMAXAREACAR 80.9288 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 406.231 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.32956 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 11.080000 0.000000 11.460000 0.700000 ;
    END
  END bot_N2MID[0]
  PIN bot_N2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.9305 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.3835 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 8.64872 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 24.7435 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.21026 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.814 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.808 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 10.5213 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 35.804 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 45.3918 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 242.56 LAYER met4  ;
    ANTENNAGATEAREA 1.3887 LAYER met4  ;
    ANTENNAMAXAREACAR 87.5954 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 453.638 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.616771 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 34.080000 0.000000 34.460000 0.700000 ;
    END
  END bot_N2END[7]
  PIN bot_N2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 19.0083 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 94.2025 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7527 LAYER met2  ;
    ANTENNAMAXAREACAR 32.3705 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 153.659 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.376412 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 11.278 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 60.616 LAYER met3  ;
    ANTENNAGATEAREA 0.7527 LAYER met3  ;
    ANTENNAMAXAREACAR 47.3539 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 234.19 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.429554 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.7996 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 15.872 LAYER met4  ;
    ANTENNAGATEAREA 1.2297 LAYER met4  ;
    ANTENNAMAXAREACAR 49.6305 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 247.098 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.490985 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 32.240000 0.000000 32.620000 0.700000 ;
    END
  END bot_N2END[6]
  PIN bot_N2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.0593 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.0275 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 9.24132 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 27.7065 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.21026 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.2509 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 9.8185 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 31.8657 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 50.9538 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 272.224 LAYER met4  ;
    ANTENNAGATEAREA 1.2297 LAYER met4  ;
    ANTENNAMAXAREACAR 69.7719 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 358.92 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.598952 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 30.860000 0.000000 31.240000 0.700000 ;
    END
  END bot_N2END[5]
  PIN bot_N2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.1911 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 30.4605 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7527 LAYER met2  ;
    ANTENNAMAXAREACAR 15.5937 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 65.3142 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.376412 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 8.7936 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 47.84 LAYER met3  ;
    ANTENNAGATEAREA 1.3887 LAYER met3  ;
    ANTENNAMAXAREACAR 41.1109 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 198.657 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.574843 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 29.480000 0.000000 29.860000 0.700000 ;
    END
  END bot_N2END[4]
  PIN bot_N2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.1699 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 25.4625 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 16.2489 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 62.473 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.21026 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 21.7595 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 116.504 LAYER met3  ;
    ANTENNAGATEAREA 0.5937 LAYER met3  ;
    ANTENNAMAXAREACAR 52.8996 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 258.707 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.709591 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 33.3282 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 179.632 LAYER met4  ;
    ANTENNAGATEAREA 1.3887 LAYER met4  ;
    ANTENNAMAXAREACAR 76.8991 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 388.059 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.967925 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 27.640000 0.000000 28.020000 0.700000 ;
    END
  END bot_N2END[3]
  PIN bot_N2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 9.3952 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 46.3925 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5937 LAYER met2  ;
    ANTENNAMAXAREACAR 28.6632 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 133.365 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.532154 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 28.2486 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 151.6 LAYER met3  ;
    ANTENNAGATEAREA 1.2297 LAYER met3  ;
    ANTENNAMAXAREACAR 51.6351 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 256.647 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 26.260000 0.000000 26.640000 0.700000 ;
    END
  END bot_N2END[2]
  PIN bot_N2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 16.3684 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 80.948 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2297 LAYER met2  ;
    ANTENNAMAXAREACAR 47.8675 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 230.321 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.46478 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 24.880000 0.000000 25.260000 0.700000 ;
    END
  END bot_N2END[1]
  PIN bot_N2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 12.3679 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 61.3445 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5937 LAYER met2  ;
    ANTENNAMAXAREACAR 25.9285 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 110.928 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.390645 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.3759 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.8 LAYER met3  ;
    ANTENNAGATEAREA 0.9117 LAYER met3  ;
    ANTENNAMAXAREACAR 30.1717 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 142.331 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.492931 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.3998 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 7.936 LAYER met4  ;
    ANTENNAGATEAREA 1.5477 LAYER met4  ;
    ANTENNAMAXAREACAR 65.1557 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 332.584 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.732075 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 23.040000 0.000000 23.420000 0.700000 ;
    END
  END bot_N2END[0]
  PIN bot_N4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.3452 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 26.565 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 103.651 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 553.744 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6312 LAYER met4  ;
    ANTENNAMAXAREACAR 181.081 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 961.837 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 58.460000 0.000000 58.840000 0.700000 ;
    END
  END bot_N4END[15]
  PIN bot_N4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1879 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.7785 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.469 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.3041 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 115.737 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 618.672 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.5006 LAYER met4  ;
    ANTENNAMAXAREACAR 87.2661 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 446.397 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 56.620000 0.000000 57.000000 0.700000 ;
    END
  END bot_N4END[14]
  PIN bot_N4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6321 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.9995 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.642 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.224 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.3041 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 118.114 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 631.824 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.5006 LAYER met4  ;
    ANTENNAMAXAREACAR 89.5172 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 458.309 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 55.240000 0.000000 55.620000 0.700000 ;
    END
  END bot_N4END[13]
  PIN bot_N4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9737 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.7075 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.988 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 21.736 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.3041 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 117.308 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 626.576 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.5006 LAYER met4  ;
    ANTENNAMAXAREACAR 102.461 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 545.276 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 53.860000 0.000000 54.240000 0.700000 ;
    END
  END bot_N4END[12]
  PIN bot_N4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7537 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.4895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.954 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 58.888 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.3041 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 113.335 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 605.392 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.5006 LAYER met4  ;
    ANTENNAMAXAREACAR 118.207 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 626.288 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 52.480000 0.000000 52.860000 0.700000 ;
    END
  END bot_N4END[11]
  PIN bot_N4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9149 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.2955 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.676 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.072 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 104.344 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 557.44 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6312 LAYER met4  ;
    ANTENNAMAXAREACAR 187.907 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 995.515 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 50.640000 0.000000 51.020000 0.700000 ;
    END
  END bot_N4END[10]
  PIN bot_N4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.5357 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.5175 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.78 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.96 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 100.882 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 538.976 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6312 LAYER met4  ;
    ANTENNAMAXAREACAR 187.249 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 990.161 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 49.260000 0.000000 49.640000 0.700000 ;
    END
  END bot_N4END[9]
  PIN bot_N4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.7251 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.4645 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.759 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 41.848 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.3041 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 115.023 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 613.92 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.5006 LAYER met4  ;
    ANTENNAMAXAREACAR 85.7021 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 437.13 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 47.880000 0.000000 48.260000 0.700000 ;
    END
  END bot_N4END[8]
  PIN bot_N4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.5421 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.3325 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 10.1256 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 31.8772 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.21026 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 16.684 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 89.448 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 48.5061 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 237.647 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 79.9704 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 427.92 LAYER met4  ;
    ANTENNAGATEAREA 1.2297 LAYER met4  ;
    ANTENNAMAXAREACAR 118.583 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 614.412 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.32956 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 46.040000 0.000000 46.420000 0.700000 ;
    END
  END bot_N4END[7]
  PIN bot_N4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.657 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.006 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 12.937 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 45.9834 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.328502 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.436 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 18.792 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 20.8413 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 89.2132 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.42052 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 96.6162 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 519.04 LAYER met4  ;
    ANTENNAGATEAREA 1.2297 LAYER met4  ;
    ANTENNAMAXAREACAR 138.235 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 715.656 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.47107 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 44.660000 0.000000 45.040000 0.700000 ;
    END
  END bot_N4END[6]
  PIN bot_N4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.9703 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.5725 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 10.8737 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 35.597 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.26202 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.2509 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 11.4509 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 39.7562 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.354037 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 79.4628 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 424.272 LAYER met4  ;
    ANTENNAGATEAREA 1.2297 LAYER met4  ;
    ANTENNAMAXAREACAR 89.8912 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 461.66 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.565409 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 43.280000 0.000000 43.660000 0.700000 ;
    END
  END bot_N4END[5]
  PIN bot_N4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.9473 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.4675 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 8.98367 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 26.4182 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.21026 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.618 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.096 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 12.7058 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 47.343 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 78.7296 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 420.832 LAYER met4  ;
    ANTENNAGATEAREA 1.2297 LAYER met4  ;
    ANTENNAMAXAREACAR 96.3728 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 500.134 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.716352 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 41.440000 0.000000 41.820000 0.700000 ;
    END
  END bot_N4END[4]
  PIN bot_N4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9737 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.7075 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.255 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 19.0641 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 103.552 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2297 LAYER met4  ;
    ANTENNAMAXAREACAR 71.2636 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 366.289 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 40.060000 0.000000 40.440000 0.700000 ;
    END
  END bot_N4END[3]
  PIN bot_N4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 17.6376 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 87.801 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5937 LAYER met2  ;
    ANTENNAMAXAREACAR 38.3003 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 172.72 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.390645 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 24.3082 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 130.576 LAYER met3  ;
    ANTENNAGATEAREA 1.0707 LAYER met3  ;
    ANTENNAMAXAREACAR 61.0034 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 294.674 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.863774 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 14.9658 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 80.288 LAYER met4  ;
    ANTENNAGATEAREA 1.2297 LAYER met4  ;
    ANTENNAMAXAREACAR 73.1737 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 359.964 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.863774 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 38.680000 0.000000 39.060000 0.700000 ;
    END
  END bot_N4END[2]
  PIN bot_N4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 20.9502 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 103.719 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2297 LAYER met2  ;
    ANTENNAMAXAREACAR 23.4171 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 98.1867 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 36.840000 0.000000 37.220000 0.700000 ;
    END
  END bot_N4END[1]
  PIN bot_N4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 11.5968 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 56.854 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2297 LAYER met2  ;
    ANTENNAMAXAREACAR 15.8907 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 72.7781 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 35.460000 0.000000 35.840000 0.700000 ;
    END
  END bot_N4END[0]
  PIN bot_NN4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6804 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.241 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.2509 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.8694 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 105.767 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 564.56 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.0659 LAYER met4  ;
    ANTENNAMAXAREACAR 152.064 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 786.849 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.820733 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 82.840000 0.000000 83.220000 0.700000 ;
    END
  END bot_NN4END[15]
  PIN bot_NN4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1445 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.5615 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.642 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.224 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.3041 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 116.405 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 621.296 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.5006 LAYER met4  ;
    ANTENNAMAXAREACAR 83.7106 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 426.985 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.31489 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 81.460000 0.000000 81.840000 0.700000 ;
    END
  END bot_NN4END[14]
  PIN bot_NN4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6321 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.9995 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.8694 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 105.926 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 566.816 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.0659 LAYER met4  ;
    ANTENNAMAXAREACAR 139.305 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 730.688 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 79.620000 0.000000 80.000000 0.700000 ;
    END
  END bot_NN4END[13]
  PIN bot_NN4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.6397 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.0375 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.987 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.064 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.3041 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 117.622 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 629.664 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.5006 LAYER met4  ;
    ANTENNAMAXAREACAR 85.4151 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 446.326 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 78.240000 0.000000 78.620000 0.700000 ;
    END
  END bot_NN4END[12]
  PIN bot_NN4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2089 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.8835 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.021 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.912 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.3041 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 116.07 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 620.448 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.5006 LAYER met4  ;
    ANTENNAMAXAREACAR 93.2804 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 478.277 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 76.860000 0.000000 77.240000 0.700000 ;
    END
  END bot_NN4END[11]
  PIN bot_NN4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6321 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.9995 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.676 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.072 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.3041 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 111.291 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 594.016 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.5006 LAYER met4  ;
    ANTENNAMAXAREACAR 103.606 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 542.744 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.706229 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 75.020000 0.000000 75.400000 0.700000 ;
    END
  END bot_NN4END[10]
  PIN bot_NN4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0667 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.1725 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.021 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.912 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.3041 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 112.936 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 603.264 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.5006 LAYER met4  ;
    ANTENNAMAXAREACAR 86.2668 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 440.427 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 73.640000 0.000000 74.020000 0.700000 ;
    END
  END bot_NN4END[9]
  PIN bot_NN4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.2623 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 21.1505 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.825 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.2 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 101.868 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 544.704 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6312 LAYER met4  ;
    ANTENNAMAXAREACAR 184.981 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 976.029 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 72.260000 0.000000 72.640000 0.700000 ;
    END
  END bot_NN4END[8]
  PIN bot_NN4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.2473 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.9675 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 7.52151 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 19.1074 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.21026 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.745 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.44 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 9.23533 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 29.3214 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 86.0256 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 459.744 LAYER met4  ;
    ANTENNAGATEAREA 0.9117 LAYER met4  ;
    ANTENNAMAXAREACAR 125.211 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 649.94 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.632495 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 70.420000 0.000000 70.800000 0.700000 ;
    END
  END bot_NN4END[7]
  PIN bot_NN4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.5245 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.3535 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 9.64067 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 29.7032 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.21026 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.884 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 15.848 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 16.2751 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 66.1606 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 86.4942 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 463.184 LAYER met4  ;
    ANTENNAGATEAREA 0.9117 LAYER met4  ;
    ANTENNAMAXAREACAR 156.993 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 831.007 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.32956 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 69.040000 0.000000 69.420000 0.700000 ;
    END
  END bot_NN4END[6]
  PIN bot_NN4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.2703 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.0725 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 8.01886 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 21.5712 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.21026 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.366 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.752 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 11.1613 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 39.4042 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 89.6085 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 478.848 LAYER met4  ;
    ANTENNAGATEAREA 0.9117 LAYER met4  ;
    ANTENNAMAXAREACAR 131.402 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 688.225 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 67.660000 0.000000 68.040000 0.700000 ;
    END
  END bot_NN4END[5]
  PIN bot_NN4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.6833 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.1375 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 16.7272 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 64.8643 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.26202 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.274 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 17.928 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 24.2588 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 106.107 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.354037 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 75.4116 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 403.136 LAYER met4  ;
    ANTENNAGATEAREA 0.7527 LAYER met4  ;
    ANTENNAMAXAREACAR 124.447 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 641.693 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.574843 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 65.820000 0.000000 66.200000 0.700000 ;
    END
  END bot_NN4END[4]
  PIN bot_NN4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7365 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.4035 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 13.1458 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 46.9577 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.26202 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.26895 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.832 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 13.7646 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 51.1721 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.354037 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 16.8375 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 90.736 LAYER met4  ;
    ANTENNAGATEAREA 0.9117 LAYER met4  ;
    ANTENNAMAXAREACAR 46.6665 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 232.17 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 64.440000 0.000000 64.820000 0.700000 ;
    END
  END bot_NN4END[3]
  PIN bot_NN4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 15.2505 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 75.7575 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5937 LAYER met2  ;
    ANTENNAMAXAREACAR 32.8193 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 145.381 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.390645 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 12.3177 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 66.16 LAYER met3  ;
    ANTENNAGATEAREA 0.9117 LAYER met3  ;
    ANTENNAMAXAREACAR 53.3881 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 263.014 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.574843 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 63.060000 0.000000 63.440000 0.700000 ;
    END
  END bot_NN4END[2]
  PIN bot_NN4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 22.4694 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 111.797 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9117 LAYER met2  ;
    ANTENNAMAXAREACAR 37.2689 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 177.452 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 61.220000 0.000000 61.600000 0.700000 ;
    END
  END bot_NN4END[1]
  PIN bot_NN4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 9.4202 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 46.403 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7527 LAYER met2  ;
    ANTENNAMAXAREACAR 19.397 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 87.089 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.46478 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 59.840000 0.000000 60.220000 0.700000 ;
    END
  END bot_NN4END[0]
  PIN UserCLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6321 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.9995 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 78.4924 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 423.672 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 10.1727 LAYER met3  ;
    ANTENNAMAXAREACAR 25.4277 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 123.135 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.578775 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.1318 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 11.84 LAYER met4  ;
    ANTENNAGATEAREA 10.4907 LAYER met4  ;
    ANTENNAMAXAREACAR 25.6309 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 124.263 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.700629 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 163.800000 0.000000 164.180000 0.700000 ;
    END
  END UserCLK
  PIN UserCLKo
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.9074 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.429 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 163.800000 399.820000 164.180000 400.520000 ;
    END
  END UserCLKo
  PIN top_FrameData[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 32.3779 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 174.08 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.5852 LAYER met3  ;
    ANTENNAMAXAREACAR 42.6731 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 213.844 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.993158 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.4388 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 40.144 LAYER met4  ;
    ANTENNAGATEAREA 2.6982 LAYER met4  ;
    ANTENNAMAXAREACAR 45.4301 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 228.722 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.993158 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 394.260000 0.700000 394.640000 ;
    END
  END top_FrameData[31]
  PIN top_FrameData[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 8.1798 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 44.552 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.6982 LAYER met3  ;
    ANTENNAMAXAREACAR 50.0168 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 245.894 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.590566 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 392.430000 0.700000 392.810000 ;
    END
  END top_FrameData[30]
  PIN top_FrameData[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 10.9468 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 58.84 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.7442 LAYER met3  ;
    ANTENNAMAXAREACAR 49.7333 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 246.138 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.482015 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 29.2977 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 156.72 LAYER met4  ;
    ANTENNAGATEAREA 2.6982 LAYER met4  ;
    ANTENNAMAXAREACAR 60.5915 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 304.221 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 391.210000 0.700000 391.590000 ;
    END
  END top_FrameData[29]
  PIN top_FrameData[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 19.793 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 107.432 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.7442 LAYER met3  ;
    ANTENNAMAXAREACAR 38.1758 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 191.153 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.872281 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 37.0785 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 198.688 LAYER met4  ;
    ANTENNAGATEAREA 2.6982 LAYER met4  ;
    ANTENNAMAXAREACAR 51.9178 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 264.79 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.872281 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 389.380000 0.700000 389.760000 ;
    END
  END top_FrameData[28]
  PIN top_FrameData[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 25.0639 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 134.136 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7527 LAYER met3  ;
    ANTENNAMAXAREACAR 53.7828 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 275.062 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.627985 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 40.4913 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 217.36 LAYER met4  ;
    ANTENNAGATEAREA 2.6982 LAYER met4  ;
    ANTENNAMAXAREACAR 76.9698 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 392.882 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.07223 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 388.160000 0.700000 388.540000 ;
    END
  END top_FrameData[27]
  PIN top_FrameData[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.7324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.368 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5937 LAYER met3  ;
    ANTENNAMAXAREACAR 18.9663 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 76.9343 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.525393 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 29.982 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 161.776 LAYER met4  ;
    ANTENNAGATEAREA 2.6982 LAYER met4  ;
    ANTENNAMAXAREACAR 58.6313 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 305.621 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.00269 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 386.330000 0.700000 386.710000 ;
    END
  END top_FrameData[26]
  PIN top_FrameData[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 23.9689 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 128.752 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.8657 LAYER met3  ;
    ANTENNAMAXAREACAR 70.621 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 351.795 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.753515 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 13.5357 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 72.656 LAYER met4  ;
    ANTENNAGATEAREA 2.6982 LAYER met4  ;
    ANTENNAMAXAREACAR 75.6376 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 378.722 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.753515 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 385.110000 0.700000 385.490000 ;
    END
  END top_FrameData[25]
  PIN top_FrameData[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 8.4925 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 46.704 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.2212 LAYER met3  ;
    ANTENNAMAXAREACAR 43.1049 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 212.24 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.592851 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 17.0268 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 91.28 LAYER met4  ;
    ANTENNAGATEAREA 2.6982 LAYER met4  ;
    ANTENNAMAXAREACAR 49.4153 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 246.07 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.674423 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 383.280000 0.700000 383.660000 ;
    END
  END top_FrameData[24]
  PIN top_FrameData[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 27.8742 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 150.984 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.5852 LAYER met3  ;
    ANTENNAMAXAREACAR 64.1385 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 323.385 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.12 LAYER via3  ;
    ANTENNAMAXCUTCAR 1.04362 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 52.5432 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 282.112 LAYER met4  ;
    ANTENNAGATEAREA 2.6982 LAYER met4  ;
    ANTENNAMAXAREACAR 83.6119 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 427.941 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04362 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 382.060000 0.700000 382.440000 ;
    END
  END top_FrameData[23]
  PIN top_FrameData[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 28.1657 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 151.136 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.0707 LAYER met3  ;
    ANTENNAMAXAREACAR 45.2115 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 231.012 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.901133 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 55.3461 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 297.056 LAYER met4  ;
    ANTENNAGATEAREA 2.6982 LAYER met4  ;
    ANTENNAMAXAREACAR 107.402 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 560.873 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.47107 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 380.840000 0.700000 381.220000 ;
    END
  END top_FrameData[22]
  PIN top_FrameData[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 17.6925 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 94.8 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9117 LAYER met3  ;
    ANTENNAMAXAREACAR 30.8017 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 142.233 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.12 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.706465 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 43.2843 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 232.256 LAYER met4  ;
    ANTENNAGATEAREA 2.6982 LAYER met4  ;
    ANTENNAMAXAREACAR 119.834 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 621.784 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 379.010000 0.700000 379.390000 ;
    END
  END top_FrameData[21]
  PIN top_FrameData[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.5044 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 19.152 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7527 LAYER met3  ;
    ANTENNAMAXAREACAR 20.6651 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 101.138 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.482697 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 34.8564 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 187.312 LAYER met4  ;
    ANTENNAGATEAREA 2.6982 LAYER met4  ;
    ANTENNAMAXAREACAR 70.5883 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 356.515 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.32956 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 377.790000 0.700000 378.170000 ;
    END
  END top_FrameData[20]
  PIN top_FrameData[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 22.548 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 120.712 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.6982 LAYER met3  ;
    ANTENNAMAXAREACAR 51.5824 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 255.892 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.574843 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 375.960000 0.700000 376.340000 ;
    END
  END top_FrameData[19]
  PIN top_FrameData[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 33.7132 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 180.736 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.7067 LAYER met3  ;
    ANTENNAMAXAREACAR 54.4901 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 274.476 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.55111 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 21.7467 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 116.448 LAYER met4  ;
    ANTENNAGATEAREA 2.6982 LAYER met4  ;
    ANTENNAMAXAREACAR 62.5498 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 317.633 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 374.740000 0.700000 375.120000 ;
    END
  END top_FrameData[18]
  PIN top_FrameData[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 12.3917 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 67 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9117 LAYER met3  ;
    ANTENNAMAXAREACAR 68.6988 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 342.747 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.870289 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.8508 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 5.008 LAYER met4  ;
    ANTENNAGATEAREA 2.6982 LAYER met4  ;
    ANTENNAMAXAREACAR 69.0141 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 344.603 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.870289 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 372.910000 0.700000 373.290000 ;
    END
  END top_FrameData[17]
  PIN top_FrameData[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 23.9775 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 128.816 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.6982 LAYER met3  ;
    ANTENNAMAXAREACAR 35.1669 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 170.806 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.590566 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 371.690000 0.700000 372.070000 ;
    END
  END top_FrameData[16]
  PIN top_FrameData[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.8034 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.08 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5937 LAYER met3  ;
    ANTENNAMAXAREACAR 25.9847 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 114.312 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.525393 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 29.5176 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 158.368 LAYER met4  ;
    ANTENNAGATEAREA 2.6982 LAYER met4  ;
    ANTENNAMAXAREACAR 58.8582 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 293.786 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.757233 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 369.860000 0.700000 370.240000 ;
    END
  END top_FrameData[15]
  PIN top_FrameData[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.1344 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 22.512 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9117 LAYER met3  ;
    ANTENNAMAXAREACAR 28.8301 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 131.405 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.596402 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 60.2964 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 326.28 LAYER met4  ;
    ANTENNAGATEAREA 2.6982 LAYER met4  ;
    ANTENNAMAXAREACAR 71.1661 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 362.574 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.967925 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 368.640000 0.700000 369.020000 ;
    END
  END top_FrameData[14]
  PIN top_FrameData[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 6.5752 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 36 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.1837 LAYER met3  ;
    ANTENNAMAXAREACAR 28.8712 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 140.635 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.539002 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 15.3723 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 83.392 LAYER met4  ;
    ANTENNAGATEAREA 2.6982 LAYER met4  ;
    ANTENNAMAXAREACAR 38.2479 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 191.181 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 367.420000 0.700000 367.800000 ;
    END
  END top_FrameData[13]
  PIN top_FrameData[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.1326 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 22.032 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 55.6161 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 298.496 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.6982 LAYER met4  ;
    ANTENNAMAXAREACAR 71.4686 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 370.936 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.32956 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 365.590000 0.700000 365.970000 ;
    END
  END top_FrameData[12]
  PIN top_FrameData[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.6634 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7527 LAYER met3  ;
    ANTENNAMAXAREACAR 17.0974 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 81.6573 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.624206 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.0676 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 11.968 LAYER met4  ;
    ANTENNAGATEAREA 2.6982 LAYER met4  ;
    ANTENNAMAXAREACAR 46.9863 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 231.089 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.624206 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 364.370000 0.700000 364.750000 ;
    END
  END top_FrameData[11]
  PIN top_FrameData[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 23.806 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 128.368 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.7067 LAYER met3  ;
    ANTENNAMAXAREACAR 47.532 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 237.836 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.797441 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.8638 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 15.744 LAYER met4  ;
    ANTENNAGATEAREA 2.6982 LAYER met4  ;
    ANTENNAMAXAREACAR 55.9006 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 280.958 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.797441 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 362.540000 0.700000 362.920000 ;
    END
  END top_FrameData[10]
  PIN top_FrameData[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 15.0431 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 80.688 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 36.7812 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 198.048 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.1045 LAYER met4  ;
    ANTENNAMAXAREACAR 56.6163 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 299.028 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 361.320000 0.700000 361.700000 ;
    END
  END top_FrameData[9]
  PIN top_FrameData[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9256 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 20.928 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 24.9297 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 133.424 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.1045 LAYER met4  ;
    ANTENNAMAXAREACAR 62.5328 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 318.273 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 359.490000 0.700000 359.870000 ;
    END
  END top_FrameData[8]
  PIN top_FrameData[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9366 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 89.9232 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 481.472 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.1045 LAYER met4  ;
    ANTENNAMAXAREACAR 106.009 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 545.93 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.920755 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 358.270000 0.700000 358.650000 ;
    END
  END top_FrameData[7]
  PIN top_FrameData[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 30.5096 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 163.176 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 13.3944 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 75.2 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.1045 LAYER met4  ;
    ANTENNAMAXAREACAR 66.6061 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 338.936 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.32956 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 356.440000 0.700000 356.820000 ;
    END
  END top_FrameData[6]
  PIN top_FrameData[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.642 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.224 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 67.4067 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 362.32 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.1045 LAYER met4  ;
    ANTENNAMAXAREACAR 82.0788 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 435.205 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.07799 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 355.220000 0.700000 355.600000 ;
    END
  END top_FrameData[5]
  PIN top_FrameData[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.2376 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 38.592 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 51.0006 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 272.944 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.1045 LAYER met4  ;
    ANTENNAMAXAREACAR 59.5482 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 305.253 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.762093 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 354.000000 0.700000 354.380000 ;
    END
  END top_FrameData[4]
  PIN top_FrameData[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 23.9856 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 130.28 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.1045 LAYER met3  ;
    ANTENNAMAXAREACAR 48.4954 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 240.516 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.967925 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 352.170000 0.700000 352.550000 ;
    END
  END top_FrameData[3]
  PIN top_FrameData[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 46.1868 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 247.728 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.113 LAYER met3  ;
    ANTENNAMAXAREACAR 70.6169 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 363.215 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.862354 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 18.7947 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 100.704 LAYER met4  ;
    ANTENNAGATEAREA 2.1045 LAYER met4  ;
    ANTENNAMAXAREACAR 79.5476 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 411.067 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.862354 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 350.950000 0.700000 351.330000 ;
    END
  END top_FrameData[2]
  PIN top_FrameData[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.6836 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 14.304 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 13.5966 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 73.456 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.1045 LAYER met4  ;
    ANTENNAMAXAREACAR 65.2225 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 332.656 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.766667 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 349.120000 0.700000 349.500000 ;
    END
  END top_FrameData[1]
  PIN top_FrameData[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.2404 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 49.744 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.636 LAYER met3  ;
    ANTENNAMAXAREACAR 59.6775 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 298.752 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.653459 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 14.5116 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 78.336 LAYER met4  ;
    ANTENNAGATEAREA 2.1045 LAYER met4  ;
    ANTENNAMAXAREACAR 66.573 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 335.975 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.737317 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 347.900000 0.700000 348.280000 ;
    END
  END top_FrameData[0]
  PIN top_FrameData_O[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 394.260000 200.100000 394.640000 ;
    END
  END top_FrameData_O[31]
  PIN top_FrameData_O[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.5404 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 13.544 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 392.430000 200.100000 392.810000 ;
    END
  END top_FrameData_O[30]
  PIN top_FrameData_O[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 391.210000 200.100000 391.590000 ;
    END
  END top_FrameData_O[29]
  PIN top_FrameData_O[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 6.4044 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 34.152 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 389.380000 200.100000 389.760000 ;
    END
  END top_FrameData_O[28]
  PIN top_FrameData_O[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 388.160000 200.100000 388.540000 ;
    END
  END top_FrameData_O[27]
  PIN top_FrameData_O[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.2614 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 12.056 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 386.330000 200.100000 386.710000 ;
    END
  END top_FrameData_O[26]
  PIN top_FrameData_O[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 385.110000 200.100000 385.490000 ;
    END
  END top_FrameData_O[25]
  PIN top_FrameData_O[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 383.280000 200.100000 383.660000 ;
    END
  END top_FrameData_O[24]
  PIN top_FrameData_O[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.5764 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 29.736 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 382.060000 200.100000 382.440000 ;
    END
  END top_FrameData_O[23]
  PIN top_FrameData_O[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 380.840000 200.100000 381.220000 ;
    END
  END top_FrameData_O[22]
  PIN top_FrameData_O[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.1604 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.184 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 379.010000 200.100000 379.390000 ;
    END
  END top_FrameData_O[21]
  PIN top_FrameData_O[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.0244 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.792 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 377.790000 200.100000 378.170000 ;
    END
  END top_FrameData_O[20]
  PIN top_FrameData_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 375.960000 200.100000 376.340000 ;
    END
  END top_FrameData_O[19]
  PIN top_FrameData_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 374.740000 200.100000 375.120000 ;
    END
  END top_FrameData_O[18]
  PIN top_FrameData_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 8.7474 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 46.648 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 372.910000 200.100000 373.290000 ;
    END
  END top_FrameData_O[17]
  PIN top_FrameData_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 371.690000 200.100000 372.070000 ;
    END
  END top_FrameData_O[16]
  PIN top_FrameData_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 369.860000 200.100000 370.240000 ;
    END
  END top_FrameData_O[15]
  PIN top_FrameData_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.4364 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.656 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 368.640000 200.100000 369.020000 ;
    END
  END top_FrameData_O[14]
  PIN top_FrameData_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 367.420000 200.100000 367.800000 ;
    END
  END top_FrameData_O[13]
  PIN top_FrameData_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.6444 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 19.432 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 365.590000 200.100000 365.970000 ;
    END
  END top_FrameData_O[12]
  PIN top_FrameData_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 364.370000 200.100000 364.750000 ;
    END
  END top_FrameData_O[11]
  PIN top_FrameData_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.7124 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.128 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 362.540000 200.100000 362.920000 ;
    END
  END top_FrameData_O[10]
  PIN top_FrameData_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 361.320000 200.100000 361.700000 ;
    END
  END top_FrameData_O[9]
  PIN top_FrameData_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.7124 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.128 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 359.490000 200.100000 359.870000 ;
    END
  END top_FrameData_O[8]
  PIN top_FrameData_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 358.270000 200.100000 358.650000 ;
    END
  END top_FrameData_O[7]
  PIN top_FrameData_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 356.440000 200.100000 356.820000 ;
    END
  END top_FrameData_O[6]
  PIN top_FrameData_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.2744 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 22.536 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 355.220000 200.100000 355.600000 ;
    END
  END top_FrameData_O[5]
  PIN top_FrameData_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.2644 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 12.072 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 354.000000 200.100000 354.380000 ;
    END
  END top_FrameData_O[4]
  PIN top_FrameData_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.7124 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.128 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 352.170000 200.100000 352.550000 ;
    END
  END top_FrameData_O[3]
  PIN top_FrameData_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 350.950000 200.100000 351.330000 ;
    END
  END top_FrameData_O[2]
  PIN top_FrameData_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.4364 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.656 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 349.120000 200.100000 349.500000 ;
    END
  END top_FrameData_O[1]
  PIN top_FrameData_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 347.900000 200.100000 348.280000 ;
    END
  END top_FrameData_O[0]
  PIN bot_FrameData[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 30.5698 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 164.912 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.5017 LAYER met3  ;
    ANTENNAMAXAREACAR 45.752 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 228.161 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.590832 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 35.3268 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 188.88 LAYER met4  ;
    ANTENNAGATEAREA 2.6982 LAYER met4  ;
    ANTENNAMAXAREACAR 58.8448 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 298.163 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 194.790000 0.700000 195.170000 ;
    END
  END bot_FrameData[31]
  PIN bot_FrameData[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 36.8044 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 197.688 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.5017 LAYER met3  ;
    ANTENNAMAXAREACAR 48.0097 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 240.137 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.983914 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 31.9608 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 170.928 LAYER met4  ;
    ANTENNAGATEAREA 2.6982 LAYER met4  ;
    ANTENNAMAXAREACAR 59.8549 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 303.486 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.983914 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 192.960000 0.700000 193.340000 ;
    END
  END bot_FrameData[30]
  PIN bot_FrameData[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 17.4514 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 93.536 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 45.5786 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 224.096 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.394295 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.8048 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 42.096 LAYER met4  ;
    ANTENNAGATEAREA 2.6982 LAYER met4  ;
    ANTENNAMAXAREACAR 49.1222 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 244.036 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.538357 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 191.740000 0.700000 192.120000 ;
    END
  END bot_FrameData[29]
  PIN bot_FrameData[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9414 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.816 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 5.4498 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 29.536 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.6982 LAYER met4  ;
    ANTENNAMAXAREACAR 55.5154 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 276.541 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.982749 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 189.910000 0.700000 190.290000 ;
    END
  END bot_FrameData[28]
  PIN bot_FrameData[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 14.3681 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 78.024 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.8657 LAYER met3  ;
    ANTENNAMAXAREACAR 54.9907 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 273.178 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.658603 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 4.8126 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 26.608 LAYER met4  ;
    ANTENNAGATEAREA 2.6982 LAYER met4  ;
    ANTENNAMAXAREACAR 56.7743 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 283.039 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 188.690000 0.700000 189.070000 ;
    END
  END bot_FrameData[27]
  PIN bot_FrameData[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.255 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5937 LAYER met3  ;
    ANTENNAMAXAREACAR 22.0301 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 92.2158 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.525393 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 19.4979 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 108.688 LAYER met4  ;
    ANTENNAGATEAREA 2.6982 LAYER met4  ;
    ANTENNAMAXAREACAR 63.7759 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 335.464 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.32956 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 186.860000 0.700000 187.240000 ;
    END
  END bot_FrameData[26]
  PIN bot_FrameData[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 31.168 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 166.696 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5937 LAYER met3  ;
    ANTENNAMAXAREACAR 62.6875 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 312.871 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.525393 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 6.5478 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 35.392 LAYER met4  ;
    ANTENNAGATEAREA 2.6982 LAYER met4  ;
    ANTENNAMAXAREACAR 65.1143 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 325.988 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.59385 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 185.640000 0.700000 186.020000 ;
    END
  END bot_FrameData[25]
  PIN bot_FrameData[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.9274 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 21.408 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5937 LAYER met3  ;
    ANTENNAMAXAREACAR 20.3794 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 79.817 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.525393 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.7996 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 15.872 LAYER met4  ;
    ANTENNAGATEAREA 2.6982 LAYER met4  ;
    ANTENNAMAXAREACAR 51.5596 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 265.684 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.80021 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 183.810000 0.700000 184.190000 ;
    END
  END bot_FrameData[24]
  PIN bot_FrameData[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 31.9287 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 171.688 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.6982 LAYER met3  ;
    ANTENNAMAXAREACAR 53.0045 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 264.91 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.574843 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 182.590000 0.700000 182.970000 ;
    END
  END bot_FrameData[23]
  PIN bot_FrameData[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 36.5547 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 195.424 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.6982 LAYER met3  ;
    ANTENNAMAXAREACAR 49.4919 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 246.896 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.571064 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 180.760000 0.700000 181.140000 ;
    END
  END bot_FrameData[22]
  PIN bot_FrameData[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 20.114 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 109.144 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.0707 LAYER met3  ;
    ANTENNAMAXAREACAR 49.8519 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 250.72 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAMAXCUTCAR 1.1527 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 24.6954 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 133.12 LAYER met4  ;
    ANTENNAGATEAREA 2.6982 LAYER met4  ;
    ANTENNAMAXAREACAR 64.7596 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 328.795 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.1527 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 179.540000 0.700000 179.920000 ;
    END
  END bot_FrameData[21]
  PIN bot_FrameData[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 21.0301 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 113.088 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.8657 LAYER met3  ;
    ANTENNAMAXAREACAR 47.2179 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 235.746 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.711586 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 27.1485 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 145.728 LAYER met4  ;
    ANTENNAGATEAREA 2.6982 LAYER met4  ;
    ANTENNAMAXAREACAR 57.2796 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 289.756 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 178.320000 0.700000 178.700000 ;
    END
  END bot_FrameData[20]
  PIN bot_FrameData[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 8.2896 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 45.152 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.6982 LAYER met4  ;
    ANTENNAMAXAREACAR 51.1923 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 257.569 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.861183 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 176.490000 0.700000 176.870000 ;
    END
  END bot_FrameData[19]
  PIN bot_FrameData[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 10.4635 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 55.792 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7527 LAYER met3  ;
    ANTENNAMAXAREACAR 22.67 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 104.734 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.429554 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 9.1197 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 49.104 LAYER met4  ;
    ANTENNAGATEAREA 2.6982 LAYER met4  ;
    ANTENNAMAXAREACAR 56.2532 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 286.591 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.602081 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 175.270000 0.700000 175.650000 ;
    END
  END bot_FrameData[18]
  PIN bot_FrameData[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 13.383 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 72.76 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.5017 LAYER met3  ;
    ANTENNAMAXAREACAR 52.8767 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 261.65 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.716618 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 13.8438 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 74.304 LAYER met4  ;
    ANTENNAGATEAREA 2.6982 LAYER met4  ;
    ANTENNAMAXAREACAR 58.0074 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 289.188 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.716618 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 173.440000 0.700000 173.820000 ;
    END
  END bot_FrameData[17]
  PIN bot_FrameData[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.32735 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 23.472 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.5392 LAYER met3  ;
    ANTENNAMAXAREACAR 41.0968 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 201.126 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.653548 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.1208 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 38.448 LAYER met4  ;
    ANTENNAGATEAREA 2.6982 LAYER met4  ;
    ANTENNAMAXAREACAR 45.268 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 226.353 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 172.220000 0.700000 172.600000 ;
    END
  END bot_FrameData[16]
  PIN bot_FrameData[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.9365 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.456 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5937 LAYER met3  ;
    ANTENNAMAXAREACAR 21.2441 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 102.779 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.734276 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 27.6138 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 150.096 LAYER met4  ;
    ANTENNAGATEAREA 2.6982 LAYER met4  ;
    ANTENNAMAXAREACAR 76.3518 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 396.04 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.32956 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 170.390000 0.700000 170.770000 ;
    END
  END bot_FrameData[15]
  PIN bot_FrameData[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 24.5939 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 131.616 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5937 LAYER met3  ;
    ANTENNAMAXAREACAR 55.4355 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 287.219 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.709591 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 59.2503 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 319.76 LAYER met4  ;
    ANTENNAGATEAREA 2.6982 LAYER met4  ;
    ANTENNAMAXAREACAR 77.3947 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 405.728 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.32956 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 169.170000 0.700000 169.550000 ;
    END
  END bot_FrameData[14]
  PIN bot_FrameData[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.2164 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 17.616 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9117 LAYER met3  ;
    ANTENNAMAXAREACAR 18.8879 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 77.4182 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.454893 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 16.0476 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 86.528 LAYER met4  ;
    ANTENNAGATEAREA 2.6982 LAYER met4  ;
    ANTENNAMAXAREACAR 61.2566 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 305.622 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.6587 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 167.340000 0.700000 167.720000 ;
    END
  END bot_FrameData[13]
  PIN bot_FrameData[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.6654 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 25.344 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 17.254 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 72.2648 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.394295 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 55.6881 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 298.88 LAYER met4  ;
    ANTENNAGATEAREA 2.6982 LAYER met4  ;
    ANTENNAMAXAREACAR 84.4295 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 435.976 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 166.120000 0.700000 166.500000 ;
    END
  END bot_FrameData[12]
  PIN bot_FrameData[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 20.968 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 112.296 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7527 LAYER met3  ;
    ANTENNAMAXAREACAR 48.2203 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 232.05 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.482697 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 39.801 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 214.144 LAYER met4  ;
    ANTENNAGATEAREA 2.6982 LAYER met4  ;
    ANTENNAMAXAREACAR 62.9713 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 311.415 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.47107 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 164.900000 0.700000 165.280000 ;
    END
  END bot_FrameData[11]
  PIN bot_FrameData[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.7324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.368 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7527 LAYER met3  ;
    ANTENNAMAXAREACAR 18.8424 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 78.2741 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.482697 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 35.1606 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 190.336 LAYER met4  ;
    ANTENNAGATEAREA 2.6982 LAYER met4  ;
    ANTENNAMAXAREACAR 46.7767 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 247.285 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 163.070000 0.700000 163.450000 ;
    END
  END bot_FrameData[10]
  PIN bot_FrameData[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 11.7938 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 63.824 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5937 LAYER met3  ;
    ANTENNAMAXAREACAR 30.9673 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 152.782 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAMAXCUTCAR 1.10267 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 26.7564 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 144.112 LAYER met4  ;
    ANTENNAGATEAREA 2.6982 LAYER met4  ;
    ANTENNAMAXAREACAR 69.0105 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 365.013 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.10267 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 161.850000 0.700000 162.230000 ;
    END
  END bot_FrameData[9]
  PIN bot_FrameData[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 20.0428 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 107.832 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.5017 LAYER met3  ;
    ANTENNAMAXAREACAR 40.575 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 200.762 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.526509 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 42.8778 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 229.152 LAYER met4  ;
    ANTENNAGATEAREA 2.6982 LAYER met4  ;
    ANTENNAMAXAREACAR 56.4662 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 285.689 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 160.020000 0.700000 160.400000 ;
    END
  END bot_FrameData[8]
  PIN bot_FrameData[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.4113 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.992 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5937 LAYER met3  ;
    ANTENNAMAXAREACAR 9.2531 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 29.0779 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.459679 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 36.0687 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 192.832 LAYER met4  ;
    ANTENNAGATEAREA 2.6982 LAYER met4  ;
    ANTENNAMAXAREACAR 97.902 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 492.145 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 158.800000 0.700000 159.180000 ;
    END
  END bot_FrameData[7]
  PIN bot_FrameData[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.7254 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.312 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5937 LAYER met3  ;
    ANTENNAMAXAREACAR 29.2023 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 141.109 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.808412 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 55.7826 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 298.448 LAYER met4  ;
    ANTENNAGATEAREA 2.6982 LAYER met4  ;
    ANTENNAMAXAREACAR 70.0496 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 356.407 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.808412 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 156.970000 0.700000 157.350000 ;
    END
  END bot_FrameData[6]
  PIN bot_FrameData[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 43.1933 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 230.808 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7527 LAYER met3  ;
    ANTENNAMAXAREACAR 72.6543 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 378.467 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.681127 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 63.3981 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 340 LAYER met4  ;
    ANTENNAGATEAREA 2.6982 LAYER met4  ;
    ANTENNAMAXAREACAR 96.1507 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 504.477 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.716352 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 155.750000 0.700000 156.130000 ;
    END
  END bot_FrameData[5]
  PIN bot_FrameData[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 35.0416 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 188.296 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.7067 LAYER met3  ;
    ANTENNAMAXAREACAR 55.5746 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 280.433 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.991362 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 45.0456 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 240.704 LAYER met4  ;
    ANTENNAGATEAREA 2.6982 LAYER met4  ;
    ANTENNAMAXAREACAR 72.2693 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 369.642 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.991362 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 153.920000 0.700000 154.300000 ;
    END
  END bot_FrameData[4]
  PIN bot_FrameData[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 24.265 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 130.816 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.3427 LAYER met3  ;
    ANTENNAMAXAREACAR 39.7567 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 197.205 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.707221 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 5.4258 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 29.408 LAYER met4  ;
    ANTENNAGATEAREA 2.6982 LAYER met4  ;
    ANTENNAMAXAREACAR 75.5574 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 394.217 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.707221 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 152.700000 0.700000 153.080000 ;
    END
  END bot_FrameData[3]
  PIN bot_FrameData[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 6.7564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 36.496 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7527 LAYER met3  ;
    ANTENNAMAXAREACAR 25.8831 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 128.583 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.482697 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 21.4356 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 117.136 LAYER met4  ;
    ANTENNAGATEAREA 2.6982 LAYER met4  ;
    ANTENNAMAXAREACAR 83.8362 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 443.639 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.32956 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 150.870000 0.700000 151.250000 ;
    END
  END bot_FrameData[2]
  PIN bot_FrameData[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 22.2226 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 119.928 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.3802 LAYER met3  ;
    ANTENNAMAXAREACAR 53.3671 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 265.613 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.665974 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 8.1066 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 44.176 LAYER met4  ;
    ANTENNAGATEAREA 2.6982 LAYER met4  ;
    ANTENNAMAXAREACAR 56.3715 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 281.986 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.665974 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 149.650000 0.700000 150.030000 ;
    END
  END bot_FrameData[1]
  PIN bot_FrameData[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.344 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 28.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 20.1444 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 108.848 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.6982 LAYER met4  ;
    ANTENNAMAXAREACAR 50.6673 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 253.34 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.32956 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 148.430000 0.700000 148.810000 ;
    END
  END bot_FrameData[0]
  PIN bot_FrameData_O[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 194.790000 200.100000 195.170000 ;
    END
  END bot_FrameData_O[31]
  PIN bot_FrameData_O[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 192.960000 200.100000 193.340000 ;
    END
  END bot_FrameData_O[30]
  PIN bot_FrameData_O[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.7124 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.128 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 191.740000 200.100000 192.120000 ;
    END
  END bot_FrameData_O[29]
  PIN bot_FrameData_O[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 189.910000 200.100000 190.290000 ;
    END
  END bot_FrameData_O[28]
  PIN bot_FrameData_O[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.7124 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.128 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 188.690000 200.100000 189.070000 ;
    END
  END bot_FrameData_O[27]
  PIN bot_FrameData_O[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 186.860000 200.100000 187.240000 ;
    END
  END bot_FrameData_O[26]
  PIN bot_FrameData_O[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.7484 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 25.32 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 185.640000 200.100000 186.020000 ;
    END
  END bot_FrameData_O[25]
  PIN bot_FrameData_O[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 183.810000 200.100000 184.190000 ;
    END
  END bot_FrameData_O[24]
  PIN bot_FrameData_O[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.9204 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 20.904 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 182.590000 200.100000 182.970000 ;
    END
  END bot_FrameData_O[23]
  PIN bot_FrameData_O[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.4244 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 23.592 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 180.760000 200.100000 181.140000 ;
    END
  END bot_FrameData_O[22]
  PIN bot_FrameData_O[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 179.540000 200.100000 179.920000 ;
    END
  END bot_FrameData_O[21]
  PIN bot_FrameData_O[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 178.320000 200.100000 178.700000 ;
    END
  END bot_FrameData_O[20]
  PIN bot_FrameData_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 176.490000 200.100000 176.870000 ;
    END
  END bot_FrameData_O[19]
  PIN bot_FrameData_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.8504 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.864 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 175.270000 200.100000 175.650000 ;
    END
  END bot_FrameData_O[18]
  PIN bot_FrameData_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 173.440000 200.100000 173.820000 ;
    END
  END bot_FrameData_O[17]
  PIN bot_FrameData_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.7124 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.128 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 172.220000 200.100000 172.600000 ;
    END
  END bot_FrameData_O[16]
  PIN bot_FrameData_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 170.390000 200.100000 170.770000 ;
    END
  END bot_FrameData_O[15]
  PIN bot_FrameData_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 169.170000 200.100000 169.550000 ;
    END
  END bot_FrameData_O[14]
  PIN bot_FrameData_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.7484 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 25.32 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 167.340000 200.100000 167.720000 ;
    END
  END bot_FrameData_O[13]
  PIN bot_FrameData_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 166.120000 200.100000 166.500000 ;
    END
  END bot_FrameData_O[12]
  PIN bot_FrameData_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 164.900000 200.100000 165.280000 ;
    END
  END bot_FrameData_O[11]
  PIN bot_FrameData_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 163.070000 200.100000 163.450000 ;
    END
  END bot_FrameData_O[10]
  PIN bot_FrameData_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.7824 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 20.168 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 161.850000 200.100000 162.230000 ;
    END
  END bot_FrameData_O[9]
  PIN bot_FrameData_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 160.020000 200.100000 160.400000 ;
    END
  END bot_FrameData_O[8]
  PIN bot_FrameData_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.8504 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.864 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 158.800000 200.100000 159.180000 ;
    END
  END bot_FrameData_O[7]
  PIN bot_FrameData_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.0694 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 27.032 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 156.970000 200.100000 157.350000 ;
    END
  END bot_FrameData_O[6]
  PIN bot_FrameData_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 155.750000 200.100000 156.130000 ;
    END
  END bot_FrameData_O[5]
  PIN bot_FrameData_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 153.920000 200.100000 154.300000 ;
    END
  END bot_FrameData_O[4]
  PIN bot_FrameData_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.7124 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.128 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 152.700000 200.100000 153.080000 ;
    END
  END bot_FrameData_O[3]
  PIN bot_FrameData_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.768 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 150.870000 200.100000 151.250000 ;
    END
  END bot_FrameData_O[2]
  PIN bot_FrameData_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 149.650000 200.100000 150.030000 ;
    END
  END bot_FrameData_O[1]
  PIN bot_FrameData_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 199.400000 148.430000 200.100000 148.810000 ;
    END
  END bot_FrameData_O[0]
  PIN FrameStrobe[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.4872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 27.426 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 36.9522 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 181.733 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.261578 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 194.160000 0.000000 194.540000 0.700000 ;
    END
  END FrameStrobe[19]
  PIN FrameStrobe[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7175 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.4265 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.538 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.336 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.8694 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 107.906 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 575.968 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.0659 LAYER met4  ;
    ANTENNAMAXAREACAR 109.951 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 567.8 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.336632 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 192.780000 0.000000 193.160000 0.700000 ;
    END
  END FrameStrobe[18]
  PIN FrameStrobe[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.2127 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.9025 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.436 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 18.792 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.8694 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 104.66 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 558.656 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.0659 LAYER met4  ;
    ANTENNAMAXAREACAR 111.422 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 573.284 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.502667 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 191.400000 0.000000 191.780000 0.700000 ;
    END
  END FrameStrobe[17]
  PIN FrameStrobe[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8883 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.2805 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.952 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.544 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.3041 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 110.063 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 587.472 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.5006 LAYER met4  ;
    ANTENNAMAXAREACAR 82.4475 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 419.149 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.31489 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 190.020000 0.000000 190.400000 0.700000 ;
    END
  END FrameStrobe[16]
  PIN FrameStrobe[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8673 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.1755 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.987 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.064 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.8694 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 108.185 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 577.456 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.0659 LAYER met4  ;
    ANTENNAMAXAREACAR 117.339 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 603.407 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.451135 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 188.180000 0.000000 188.560000 0.700000 ;
    END
  END FrameStrobe[15]
  PIN FrameStrobe[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 19.6107 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 95.0254 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.261578 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 186.800000 0.000000 187.180000 0.700000 ;
    END
  END FrameStrobe[14]
  PIN FrameStrobe[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2512 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.246 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 23.1201 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 108.934 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.261578 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 185.420000 0.000000 185.800000 0.700000 ;
    END
  END FrameStrobe[13]
  PIN FrameStrobe[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6321 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.9995 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.255 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 47.0856 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 252.064 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.7192 LAYER met4  ;
    ANTENNAMAXAREACAR 50.5547 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 246.963 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.695197 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 183.580000 0.000000 183.960000 0.700000 ;
    END
  END FrameStrobe[12]
  PIN FrameStrobe[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 47.7569 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 236.688 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.4557 LAYER met2  ;
    ANTENNAMAXAREACAR 35.9703 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 169.661 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.476355 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.5798 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 24.896 LAYER met3  ;
    ANTENNAGATEAREA 5.7192 LAYER met3  ;
    ANTENNAMAXAREACAR 36.771 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 174.014 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.482452 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 182.200000 0.000000 182.580000 0.700000 ;
    END
  END FrameStrobe[11]
  PIN FrameStrobe[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 31.289 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 154.21 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.8112 LAYER met2  ;
    ANTENNAMAXAREACAR 34.4437 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 165.969 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.616785 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 9.8628 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 53.072 LAYER met3  ;
    ANTENNAGATEAREA 5.7192 LAYER met3  ;
    ANTENNAMAXAREACAR 36.1682 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 175.248 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.616785 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 180.820000 0.000000 181.200000 0.700000 ;
    END
  END FrameStrobe[10]
  PIN FrameStrobe[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8029 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.8535 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 20.824 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 111.528 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 21.0192 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 113.984 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.7192 LAYER met4  ;
    ANTENNAMAXAREACAR 37.2664 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 187.864 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.967925 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 178.980000 0.000000 179.360000 0.700000 ;
    END
  END FrameStrobe[9]
  PIN FrameStrobe[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.2473 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.9675 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 7.52151 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 19.1074 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.21026 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 9.301 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 50.072 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 28.9179 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 134.295 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 13.8438 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 74.304 LAYER met4  ;
    ANTENNAGATEAREA 5.7192 LAYER met4  ;
    ANTENNAMAXAREACAR 31.3385 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 147.287 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.590925 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 177.600000 0.000000 177.980000 0.700000 ;
    END
  END FrameStrobe[8]
  PIN FrameStrobe[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.0347 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.8945 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met2  ;
    ANTENNAMAXAREACAR 9.366 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 28.2137 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.26202 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 10.2862 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 34.1948 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.354037 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 30.5448 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 163.376 LAYER met4  ;
    ANTENNAGATEAREA 5.7192 LAYER met4  ;
    ANTENNAMAXAREACAR 33.7836 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 162.183 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.632332 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 176.220000 0.000000 176.600000 0.700000 ;
    END
  END FrameStrobe[7]
  PIN FrameStrobe[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6321 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.9995 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.255 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 43.5315 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 233.104 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.7192 LAYER met4  ;
    ANTENNAMAXAREACAR 28.2314 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 138.769 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.511053 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 174.380000 0.000000 174.760000 0.700000 ;
    END
  END FrameStrobe[6]
  PIN FrameStrobe[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.8921 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.2995 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 6.7479 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 36.432 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4347 LAYER met3  ;
    ANTENNAMAXAREACAR 20.3812 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 89.8252 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.302277 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 32.6364 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 175.472 LAYER met4  ;
    ANTENNAGATEAREA 5.7192 LAYER met4  ;
    ANTENNAMAXAREACAR 36.2826 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 173.522 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.658603 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 173.000000 0.000000 173.380000 0.700000 ;
    END
  END FrameStrobe[5]
  PIN FrameStrobe[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 15.1371 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 74.1685 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.7067 LAYER met2  ;
    ANTENNAMAXAREACAR 21.3224 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 101.11 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.488217 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.815 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 15.48 LAYER met3  ;
    ANTENNAGATEAREA 1.7067 LAYER met3  ;
    ANTENNAMAXAREACAR 22.9717 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 110.18 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.511654 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 50.0532 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 268.832 LAYER met4  ;
    ANTENNAGATEAREA 5.7192 LAYER met4  ;
    ANTENNAMAXAREACAR 66.958 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 350.368 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.47107 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 171.620000 0.000000 172.000000 0.700000 ;
    END
  END FrameStrobe[4]
  PIN FrameStrobe[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 23.3763 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 114.86 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.3427 LAYER met2  ;
    ANTENNAMAXAREACAR 22.7683 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 108.673 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.781947 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 8.4538 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 46.024 LAYER met3  ;
    ANTENNAGATEAREA 4.2507 LAYER met3  ;
    ANTENNAMAXAREACAR 24.7571 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 119.501 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.791358 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 22.0626 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 118.608 LAYER met4  ;
    ANTENNAGATEAREA 5.7192 LAYER met4  ;
    ANTENNAMAXAREACAR 55.0236 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 282.696 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.798482 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 169.780000 0.000000 170.160000 0.700000 ;
    END
  END FrameStrobe[3]
  PIN FrameStrobe[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.1788 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 65.065 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3887 LAYER met2  ;
    ANTENNAMAXAREACAR 17.8956 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 81.2274 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.493584 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 34.3434 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 184.576 LAYER met3  ;
    ANTENNAGATEAREA 5.7192 LAYER met3  ;
    ANTENNAMAXAREACAR 35.5101 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 170.041 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.527673 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 168.400000 0.000000 168.780000 0.700000 ;
    END
  END FrameStrobe[2]
  PIN FrameStrobe[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 11.4796 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 56.343 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.7067 LAYER met2  ;
    ANTENNAMAXAREACAR 22.2463 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 101.214 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.488217 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 16.2508 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 87.608 LAYER met3  ;
    ANTENNAGATEAREA 2.3427 LAYER met3  ;
    ANTENNAMAXAREACAR 29.1831 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 138.61 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.505291 LAYER via3  ;
    ANTENNADIFFAREA 0.4347 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 15.2916 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 82.496 LAYER met4  ;
    ANTENNAGATEAREA 5.7192 LAYER met4  ;
    ANTENNAMAXAREACAR 36.0193 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 179.975 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.569602 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 167.020000 0.000000 167.400000 0.700000 ;
    END
  END FrameStrobe[1]
  PIN FrameStrobe[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 38.4588 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 188.482 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.7192 LAYER met2  ;
    ANTENNAMAXAREACAR 21.8654 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 104.355 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.523155 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 165.180000 0.000000 165.560000 0.700000 ;
    END
  END FrameStrobe[0]
  PIN FrameStrobe_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.3998 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.891 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 194.160000 399.820000 194.540000 400.520000 ;
    END
  END FrameStrobe_O[19]
  PIN FrameStrobe_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.8586 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 24.185 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 192.780000 399.820000 193.160000 400.520000 ;
    END
  END FrameStrobe_O[18]
  PIN FrameStrobe_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.511 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 27.447 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 191.400000 399.820000 191.780000 400.520000 ;
    END
  END FrameStrobe_O[17]
  PIN FrameStrobe_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.8926 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.355 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 190.020000 399.820000 190.400000 400.520000 ;
    END
  END FrameStrobe_O[16]
  PIN FrameStrobe_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.531 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 22.547 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 188.180000 399.820000 188.560000 400.520000 ;
    END
  END FrameStrobe_O[15]
  PIN FrameStrobe_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.283 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 21.189 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 186.800000 399.820000 187.180000 400.520000 ;
    END
  END FrameStrobe_O[14]
  PIN FrameStrobe_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.019 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.987 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 185.420000 399.820000 185.800000 400.520000 ;
    END
  END FrameStrobe_O[13]
  PIN FrameStrobe_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.4146 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.965 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 183.580000 399.820000 183.960000 400.520000 ;
    END
  END FrameStrobe_O[12]
  PIN FrameStrobe_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.8122 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.953 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 182.200000 399.820000 182.580000 400.520000 ;
    END
  END FrameStrobe_O[11]
  PIN FrameStrobe_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.6386 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.085 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 180.820000 399.820000 181.200000 400.520000 ;
    END
  END FrameStrobe_O[10]
  PIN FrameStrobe_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.1782 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 20.783 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 178.980000 399.820000 179.360000 400.520000 ;
    END
  END FrameStrobe_O[9]
  PIN FrameStrobe_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.3694 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.739 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 177.600000 399.820000 177.980000 400.520000 ;
    END
  END FrameStrobe_O[8]
  PIN FrameStrobe_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.8926 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.355 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 176.220000 399.820000 176.600000 400.520000 ;
    END
  END FrameStrobe_O[7]
  PIN FrameStrobe_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.3662 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.723 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 174.380000 399.820000 174.760000 400.520000 ;
    END
  END FrameStrobe_O[6]
  PIN FrameStrobe_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0437 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.0575 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.7968 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 20.72 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 173.000000 399.820000 173.380000 400.520000 ;
    END
  END FrameStrobe_O[5]
  PIN FrameStrobe_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.479 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.287 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 171.620000 399.820000 172.000000 400.520000 ;
    END
  END FrameStrobe_O[4]
  PIN FrameStrobe_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.1458 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.621 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 169.780000 399.820000 170.160000 400.520000 ;
    END
  END FrameStrobe_O[3]
  PIN FrameStrobe_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.0506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.145 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 168.400000 399.820000 168.780000 400.520000 ;
    END
  END FrameStrobe_O[2]
  PIN FrameStrobe_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.1078 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.313 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 167.020000 399.820000 167.400000 400.520000 ;
    END
  END FrameStrobe_O[1]
  PIN FrameStrobe_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.305 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.417 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 165.180000 399.820000 165.560000 400.520000 ;
    END
  END FrameStrobe_O[0]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 198.900000 395.790000 200.100000 396.990000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000000 395.790000 1.200000 396.990000 ;
    END
    PORT
      LAYER met3 ;
        RECT 198.900000 2.850000 200.100000 4.050000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000000 2.850000 1.200000 4.050000 ;
    END
    PORT
      LAYER met4 ;
        RECT 196.070000 399.320000 197.270000 400.520000 ;
    END
    PORT
      LAYER met4 ;
        RECT 196.070000 0.000000 197.270000 1.200000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2.830000 399.320000 4.030000 400.520000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2.830000 0.000000 4.030000 1.200000 ;
    END

# P/G power stripe data as pin
    PORT
      LAYER met3 ;
        RECT 0.000000 2.850000 200.100000 4.050000 ;
        RECT 0.000000 395.790000 200.100000 396.990000 ;
        RECT 2.830000 4.860000 4.030000 5.340000 ;
        RECT 2.830000 10.300000 4.030000 10.780000 ;
        RECT 7.060000 4.860000 8.260000 5.340000 ;
        RECT 7.060000 10.300000 8.260000 10.780000 ;
        RECT 2.830000 15.740000 4.030000 16.220000 ;
        RECT 7.060000 15.740000 8.260000 16.220000 ;
        RECT 2.830000 21.180000 4.030000 21.660000 ;
        RECT 7.060000 21.180000 8.260000 21.660000 ;
        RECT 2.830000 37.500000 4.030000 37.980000 ;
        RECT 7.060000 37.500000 8.260000 37.980000 ;
        RECT 2.830000 26.620000 4.030000 27.100000 ;
        RECT 7.060000 26.620000 8.260000 27.100000 ;
        RECT 2.830000 32.060000 4.030000 32.540000 ;
        RECT 7.060000 32.060000 8.260000 32.540000 ;
        RECT 2.830000 42.940000 4.030000 43.420000 ;
        RECT 7.060000 42.940000 8.260000 43.420000 ;
        RECT 2.830000 48.380000 4.030000 48.860000 ;
        RECT 7.060000 48.380000 8.260000 48.860000 ;
        RECT 52.060000 21.180000 53.260000 21.660000 ;
        RECT 52.060000 15.740000 53.260000 16.220000 ;
        RECT 52.060000 10.300000 53.260000 10.780000 ;
        RECT 52.060000 4.860000 53.260000 5.340000 ;
        RECT 97.060000 21.180000 98.260000 21.660000 ;
        RECT 97.060000 15.740000 98.260000 16.220000 ;
        RECT 97.060000 10.300000 98.260000 10.780000 ;
        RECT 97.060000 4.860000 98.260000 5.340000 ;
        RECT 52.060000 26.620000 53.260000 27.100000 ;
        RECT 52.060000 32.060000 53.260000 32.540000 ;
        RECT 52.060000 37.500000 53.260000 37.980000 ;
        RECT 52.060000 42.940000 53.260000 43.420000 ;
        RECT 52.060000 48.380000 53.260000 48.860000 ;
        RECT 97.060000 26.620000 98.260000 27.100000 ;
        RECT 97.060000 32.060000 98.260000 32.540000 ;
        RECT 97.060000 37.500000 98.260000 37.980000 ;
        RECT 97.060000 42.940000 98.260000 43.420000 ;
        RECT 97.060000 48.380000 98.260000 48.860000 ;
        RECT 2.830000 53.820000 4.030000 54.300000 ;
        RECT 7.060000 53.820000 8.260000 54.300000 ;
        RECT 2.830000 59.260000 4.030000 59.740000 ;
        RECT 7.060000 59.260000 8.260000 59.740000 ;
        RECT 2.830000 64.700000 4.030000 65.180000 ;
        RECT 7.060000 64.700000 8.260000 65.180000 ;
        RECT 2.830000 70.140000 4.030000 70.620000 ;
        RECT 7.060000 70.140000 8.260000 70.620000 ;
        RECT 7.060000 81.020000 8.260000 81.500000 ;
        RECT 2.830000 81.020000 4.030000 81.500000 ;
        RECT 2.830000 75.580000 4.030000 76.060000 ;
        RECT 7.060000 75.580000 8.260000 76.060000 ;
        RECT 2.830000 86.460000 4.030000 86.940000 ;
        RECT 7.060000 86.460000 8.260000 86.940000 ;
        RECT 2.830000 91.900000 4.030000 92.380000 ;
        RECT 7.060000 91.900000 8.260000 92.380000 ;
        RECT 2.830000 97.340000 4.030000 97.820000 ;
        RECT 7.060000 97.340000 8.260000 97.820000 ;
        RECT 52.060000 70.140000 53.260000 70.620000 ;
        RECT 52.060000 53.820000 53.260000 54.300000 ;
        RECT 52.060000 59.260000 53.260000 59.740000 ;
        RECT 52.060000 64.700000 53.260000 65.180000 ;
        RECT 97.060000 53.820000 98.260000 54.300000 ;
        RECT 97.060000 59.260000 98.260000 59.740000 ;
        RECT 97.060000 64.700000 98.260000 65.180000 ;
        RECT 97.060000 70.140000 98.260000 70.620000 ;
        RECT 52.060000 75.580000 53.260000 76.060000 ;
        RECT 52.060000 81.020000 53.260000 81.500000 ;
        RECT 52.060000 86.460000 53.260000 86.940000 ;
        RECT 52.060000 91.900000 53.260000 92.380000 ;
        RECT 52.060000 97.340000 53.260000 97.820000 ;
        RECT 97.060000 75.580000 98.260000 76.060000 ;
        RECT 97.060000 81.020000 98.260000 81.500000 ;
        RECT 97.060000 86.460000 98.260000 86.940000 ;
        RECT 97.060000 91.900000 98.260000 92.380000 ;
        RECT 97.060000 97.340000 98.260000 97.820000 ;
        RECT 2.830000 102.780000 4.030000 103.260000 ;
        RECT 7.060000 102.780000 8.260000 103.260000 ;
        RECT 2.830000 108.220000 4.030000 108.700000 ;
        RECT 7.060000 108.220000 8.260000 108.700000 ;
        RECT 2.830000 113.660000 4.030000 114.140000 ;
        RECT 7.060000 113.660000 8.260000 114.140000 ;
        RECT 2.830000 119.100000 4.030000 119.580000 ;
        RECT 2.830000 124.540000 4.030000 125.020000 ;
        RECT 7.060000 119.100000 8.260000 119.580000 ;
        RECT 7.060000 124.540000 8.260000 125.020000 ;
        RECT 2.830000 129.980000 4.030000 130.460000 ;
        RECT 7.060000 129.980000 8.260000 130.460000 ;
        RECT 2.830000 135.420000 4.030000 135.900000 ;
        RECT 7.060000 135.420000 8.260000 135.900000 ;
        RECT 2.830000 140.860000 4.030000 141.340000 ;
        RECT 7.060000 140.860000 8.260000 141.340000 ;
        RECT 2.830000 146.300000 4.030000 146.780000 ;
        RECT 7.060000 146.300000 8.260000 146.780000 ;
        RECT 52.060000 124.540000 53.260000 125.020000 ;
        RECT 52.060000 119.100000 53.260000 119.580000 ;
        RECT 52.060000 102.780000 53.260000 103.260000 ;
        RECT 52.060000 108.220000 53.260000 108.700000 ;
        RECT 52.060000 113.660000 53.260000 114.140000 ;
        RECT 97.060000 124.540000 98.260000 125.020000 ;
        RECT 97.060000 102.780000 98.260000 103.260000 ;
        RECT 97.060000 108.220000 98.260000 108.700000 ;
        RECT 97.060000 113.660000 98.260000 114.140000 ;
        RECT 97.060000 119.100000 98.260000 119.580000 ;
        RECT 52.060000 129.980000 53.260000 130.460000 ;
        RECT 52.060000 135.420000 53.260000 135.900000 ;
        RECT 52.060000 140.860000 53.260000 141.340000 ;
        RECT 52.060000 146.300000 53.260000 146.780000 ;
        RECT 97.060000 129.980000 98.260000 130.460000 ;
        RECT 97.060000 135.420000 98.260000 135.900000 ;
        RECT 97.060000 140.860000 98.260000 141.340000 ;
        RECT 97.060000 146.300000 98.260000 146.780000 ;
        RECT 2.830000 162.620000 4.030000 163.100000 ;
        RECT 7.060000 162.620000 8.260000 163.100000 ;
        RECT 2.830000 151.740000 4.030000 152.220000 ;
        RECT 7.060000 151.740000 8.260000 152.220000 ;
        RECT 2.830000 157.180000 4.030000 157.660000 ;
        RECT 7.060000 157.180000 8.260000 157.660000 ;
        RECT 2.830000 168.060000 4.030000 168.540000 ;
        RECT 7.060000 168.060000 8.260000 168.540000 ;
        RECT 2.830000 173.500000 4.030000 173.980000 ;
        RECT 7.060000 173.500000 8.260000 173.980000 ;
        RECT 2.830000 178.940000 4.030000 179.420000 ;
        RECT 7.060000 178.940000 8.260000 179.420000 ;
        RECT 2.830000 184.380000 4.030000 184.860000 ;
        RECT 7.060000 184.380000 8.260000 184.860000 ;
        RECT 2.830000 189.820000 4.030000 190.300000 ;
        RECT 7.060000 189.820000 8.260000 190.300000 ;
        RECT 2.830000 195.260000 4.030000 195.740000 ;
        RECT 7.060000 195.260000 8.260000 195.740000 ;
        RECT 52.060000 173.500000 53.260000 173.980000 ;
        RECT 52.060000 168.060000 53.260000 168.540000 ;
        RECT 52.060000 151.740000 53.260000 152.220000 ;
        RECT 52.060000 157.180000 53.260000 157.660000 ;
        RECT 52.060000 162.620000 53.260000 163.100000 ;
        RECT 97.060000 173.500000 98.260000 173.980000 ;
        RECT 97.060000 151.740000 98.260000 152.220000 ;
        RECT 97.060000 157.180000 98.260000 157.660000 ;
        RECT 97.060000 162.620000 98.260000 163.100000 ;
        RECT 97.060000 168.060000 98.260000 168.540000 ;
        RECT 52.060000 178.940000 53.260000 179.420000 ;
        RECT 52.060000 184.380000 53.260000 184.860000 ;
        RECT 52.060000 189.820000 53.260000 190.300000 ;
        RECT 52.060000 195.260000 53.260000 195.740000 ;
        RECT 97.060000 178.940000 98.260000 179.420000 ;
        RECT 97.060000 184.380000 98.260000 184.860000 ;
        RECT 97.060000 189.820000 98.260000 190.300000 ;
        RECT 97.060000 195.260000 98.260000 195.740000 ;
        RECT 142.060000 4.860000 143.260000 5.340000 ;
        RECT 142.060000 10.300000 143.260000 10.780000 ;
        RECT 142.060000 15.740000 143.260000 16.220000 ;
        RECT 142.060000 21.180000 143.260000 21.660000 ;
        RECT 142.060000 26.620000 143.260000 27.100000 ;
        RECT 142.060000 32.060000 143.260000 32.540000 ;
        RECT 142.060000 37.500000 143.260000 37.980000 ;
        RECT 142.060000 42.940000 143.260000 43.420000 ;
        RECT 142.060000 48.380000 143.260000 48.860000 ;
        RECT 196.070000 4.860000 197.270000 5.340000 ;
        RECT 196.070000 10.300000 197.270000 10.780000 ;
        RECT 187.060000 4.860000 188.260000 5.340000 ;
        RECT 187.060000 10.300000 188.260000 10.780000 ;
        RECT 187.060000 15.740000 188.260000 16.220000 ;
        RECT 187.060000 21.180000 188.260000 21.660000 ;
        RECT 196.070000 21.180000 197.270000 21.660000 ;
        RECT 196.070000 15.740000 197.270000 16.220000 ;
        RECT 196.070000 37.500000 197.270000 37.980000 ;
        RECT 187.060000 37.500000 188.260000 37.980000 ;
        RECT 196.070000 26.620000 197.270000 27.100000 ;
        RECT 196.070000 32.060000 197.270000 32.540000 ;
        RECT 187.060000 26.620000 188.260000 27.100000 ;
        RECT 187.060000 32.060000 188.260000 32.540000 ;
        RECT 196.070000 42.940000 197.270000 43.420000 ;
        RECT 196.070000 48.380000 197.270000 48.860000 ;
        RECT 187.060000 42.940000 188.260000 43.420000 ;
        RECT 187.060000 48.380000 188.260000 48.860000 ;
        RECT 142.060000 70.140000 143.260000 70.620000 ;
        RECT 142.060000 64.700000 143.260000 65.180000 ;
        RECT 142.060000 59.260000 143.260000 59.740000 ;
        RECT 142.060000 53.820000 143.260000 54.300000 ;
        RECT 142.060000 75.580000 143.260000 76.060000 ;
        RECT 142.060000 81.020000 143.260000 81.500000 ;
        RECT 142.060000 86.460000 143.260000 86.940000 ;
        RECT 142.060000 91.900000 143.260000 92.380000 ;
        RECT 142.060000 97.340000 143.260000 97.820000 ;
        RECT 187.060000 59.260000 188.260000 59.740000 ;
        RECT 187.060000 53.820000 188.260000 54.300000 ;
        RECT 196.070000 59.260000 197.270000 59.740000 ;
        RECT 196.070000 53.820000 197.270000 54.300000 ;
        RECT 196.070000 64.700000 197.270000 65.180000 ;
        RECT 196.070000 70.140000 197.270000 70.620000 ;
        RECT 187.060000 70.140000 188.260000 70.620000 ;
        RECT 187.060000 64.700000 188.260000 65.180000 ;
        RECT 187.060000 75.580000 188.260000 76.060000 ;
        RECT 187.060000 81.020000 188.260000 81.500000 ;
        RECT 187.060000 86.460000 188.260000 86.940000 ;
        RECT 196.070000 86.460000 197.270000 86.940000 ;
        RECT 196.070000 81.020000 197.270000 81.500000 ;
        RECT 196.070000 75.580000 197.270000 76.060000 ;
        RECT 196.070000 91.900000 197.270000 92.380000 ;
        RECT 196.070000 97.340000 197.270000 97.820000 ;
        RECT 187.060000 91.900000 188.260000 92.380000 ;
        RECT 187.060000 97.340000 188.260000 97.820000 ;
        RECT 142.060000 124.540000 143.260000 125.020000 ;
        RECT 142.060000 119.100000 143.260000 119.580000 ;
        RECT 142.060000 113.660000 143.260000 114.140000 ;
        RECT 142.060000 108.220000 143.260000 108.700000 ;
        RECT 142.060000 102.780000 143.260000 103.260000 ;
        RECT 142.060000 129.980000 143.260000 130.460000 ;
        RECT 142.060000 135.420000 143.260000 135.900000 ;
        RECT 142.060000 140.860000 143.260000 141.340000 ;
        RECT 142.060000 146.300000 143.260000 146.780000 ;
        RECT 196.070000 102.780000 197.270000 103.260000 ;
        RECT 196.070000 108.220000 197.270000 108.700000 ;
        RECT 187.060000 108.220000 188.260000 108.700000 ;
        RECT 187.060000 102.780000 188.260000 103.260000 ;
        RECT 187.060000 124.540000 188.260000 125.020000 ;
        RECT 187.060000 119.100000 188.260000 119.580000 ;
        RECT 187.060000 113.660000 188.260000 114.140000 ;
        RECT 196.070000 124.540000 197.270000 125.020000 ;
        RECT 196.070000 119.100000 197.270000 119.580000 ;
        RECT 196.070000 113.660000 197.270000 114.140000 ;
        RECT 196.070000 129.980000 197.270000 130.460000 ;
        RECT 196.070000 135.420000 197.270000 135.900000 ;
        RECT 187.060000 129.980000 188.260000 130.460000 ;
        RECT 187.060000 135.420000 188.260000 135.900000 ;
        RECT 187.060000 140.860000 188.260000 141.340000 ;
        RECT 187.060000 146.300000 188.260000 146.780000 ;
        RECT 196.070000 146.300000 197.270000 146.780000 ;
        RECT 196.070000 140.860000 197.270000 141.340000 ;
        RECT 142.060000 173.500000 143.260000 173.980000 ;
        RECT 142.060000 168.060000 143.260000 168.540000 ;
        RECT 142.060000 162.620000 143.260000 163.100000 ;
        RECT 142.060000 157.180000 143.260000 157.660000 ;
        RECT 142.060000 151.740000 143.260000 152.220000 ;
        RECT 142.060000 178.940000 143.260000 179.420000 ;
        RECT 142.060000 184.380000 143.260000 184.860000 ;
        RECT 142.060000 189.820000 143.260000 190.300000 ;
        RECT 142.060000 195.260000 143.260000 195.740000 ;
        RECT 196.070000 162.620000 197.270000 163.100000 ;
        RECT 187.060000 162.620000 188.260000 163.100000 ;
        RECT 196.070000 151.740000 197.270000 152.220000 ;
        RECT 196.070000 157.180000 197.270000 157.660000 ;
        RECT 187.060000 157.180000 188.260000 157.660000 ;
        RECT 187.060000 151.740000 188.260000 152.220000 ;
        RECT 196.070000 168.060000 197.270000 168.540000 ;
        RECT 196.070000 173.500000 197.270000 173.980000 ;
        RECT 187.060000 173.500000 188.260000 173.980000 ;
        RECT 187.060000 168.060000 188.260000 168.540000 ;
        RECT 187.060000 178.940000 188.260000 179.420000 ;
        RECT 187.060000 184.380000 188.260000 184.860000 ;
        RECT 196.070000 184.380000 197.270000 184.860000 ;
        RECT 196.070000 178.940000 197.270000 179.420000 ;
        RECT 196.070000 189.820000 197.270000 190.300000 ;
        RECT 196.070000 195.260000 197.270000 195.740000 ;
        RECT 187.060000 189.820000 188.260000 190.300000 ;
        RECT 187.060000 195.260000 188.260000 195.740000 ;
        RECT 7.060000 206.140000 8.260000 206.620000 ;
        RECT 2.830000 206.140000 4.030000 206.620000 ;
        RECT 2.830000 200.700000 4.030000 201.180000 ;
        RECT 7.060000 200.700000 8.260000 201.180000 ;
        RECT 2.830000 211.580000 4.030000 212.060000 ;
        RECT 7.060000 211.580000 8.260000 212.060000 ;
        RECT 2.830000 217.020000 4.030000 217.500000 ;
        RECT 7.060000 217.020000 8.260000 217.500000 ;
        RECT 2.830000 222.460000 4.030000 222.940000 ;
        RECT 7.060000 222.460000 8.260000 222.940000 ;
        RECT 2.830000 227.900000 4.030000 228.380000 ;
        RECT 7.060000 227.900000 8.260000 228.380000 ;
        RECT 2.830000 233.340000 4.030000 233.820000 ;
        RECT 7.060000 233.340000 8.260000 233.820000 ;
        RECT 2.830000 238.780000 4.030000 239.260000 ;
        RECT 7.060000 238.780000 8.260000 239.260000 ;
        RECT 2.830000 244.220000 4.030000 244.700000 ;
        RECT 2.830000 249.660000 4.030000 250.140000 ;
        RECT 7.060000 244.220000 8.260000 244.700000 ;
        RECT 7.060000 249.660000 8.260000 250.140000 ;
        RECT 52.060000 222.460000 53.260000 222.940000 ;
        RECT 52.060000 217.020000 53.260000 217.500000 ;
        RECT 52.060000 211.580000 53.260000 212.060000 ;
        RECT 52.060000 206.140000 53.260000 206.620000 ;
        RECT 52.060000 200.700000 53.260000 201.180000 ;
        RECT 97.060000 222.460000 98.260000 222.940000 ;
        RECT 97.060000 211.580000 98.260000 212.060000 ;
        RECT 97.060000 206.140000 98.260000 206.620000 ;
        RECT 97.060000 200.700000 98.260000 201.180000 ;
        RECT 97.060000 217.020000 98.260000 217.500000 ;
        RECT 52.060000 227.900000 53.260000 228.380000 ;
        RECT 52.060000 233.340000 53.260000 233.820000 ;
        RECT 52.060000 238.780000 53.260000 239.260000 ;
        RECT 52.060000 244.220000 53.260000 244.700000 ;
        RECT 52.060000 249.660000 53.260000 250.140000 ;
        RECT 97.060000 227.900000 98.260000 228.380000 ;
        RECT 97.060000 233.340000 98.260000 233.820000 ;
        RECT 97.060000 238.780000 98.260000 239.260000 ;
        RECT 97.060000 244.220000 98.260000 244.700000 ;
        RECT 97.060000 249.660000 98.260000 250.140000 ;
        RECT 2.830000 255.100000 4.030000 255.580000 ;
        RECT 7.060000 255.100000 8.260000 255.580000 ;
        RECT 2.830000 260.540000 4.030000 261.020000 ;
        RECT 7.060000 260.540000 8.260000 261.020000 ;
        RECT 2.830000 265.980000 4.030000 266.460000 ;
        RECT 7.060000 265.980000 8.260000 266.460000 ;
        RECT 2.830000 271.420000 4.030000 271.900000 ;
        RECT 7.060000 271.420000 8.260000 271.900000 ;
        RECT 2.830000 287.740000 4.030000 288.220000 ;
        RECT 7.060000 287.740000 8.260000 288.220000 ;
        RECT 2.830000 276.860000 4.030000 277.340000 ;
        RECT 7.060000 276.860000 8.260000 277.340000 ;
        RECT 2.830000 282.300000 4.030000 282.780000 ;
        RECT 7.060000 282.300000 8.260000 282.780000 ;
        RECT 2.830000 293.180000 4.030000 293.660000 ;
        RECT 7.060000 293.180000 8.260000 293.660000 ;
        RECT 2.830000 298.620000 4.030000 299.100000 ;
        RECT 7.060000 298.620000 8.260000 299.100000 ;
        RECT 52.060000 271.420000 53.260000 271.900000 ;
        RECT 52.060000 255.100000 53.260000 255.580000 ;
        RECT 52.060000 260.540000 53.260000 261.020000 ;
        RECT 52.060000 265.980000 53.260000 266.460000 ;
        RECT 97.060000 255.100000 98.260000 255.580000 ;
        RECT 97.060000 260.540000 98.260000 261.020000 ;
        RECT 97.060000 265.980000 98.260000 266.460000 ;
        RECT 97.060000 271.420000 98.260000 271.900000 ;
        RECT 52.060000 276.860000 53.260000 277.340000 ;
        RECT 52.060000 282.300000 53.260000 282.780000 ;
        RECT 52.060000 287.740000 53.260000 288.220000 ;
        RECT 52.060000 293.180000 53.260000 293.660000 ;
        RECT 52.060000 298.620000 53.260000 299.100000 ;
        RECT 97.060000 276.860000 98.260000 277.340000 ;
        RECT 97.060000 282.300000 98.260000 282.780000 ;
        RECT 97.060000 287.740000 98.260000 288.220000 ;
        RECT 97.060000 293.180000 98.260000 293.660000 ;
        RECT 97.060000 298.620000 98.260000 299.100000 ;
        RECT 2.830000 304.060000 4.030000 304.540000 ;
        RECT 7.060000 304.060000 8.260000 304.540000 ;
        RECT 2.830000 309.500000 4.030000 309.980000 ;
        RECT 7.060000 309.500000 8.260000 309.980000 ;
        RECT 2.830000 314.940000 4.030000 315.420000 ;
        RECT 7.060000 314.940000 8.260000 315.420000 ;
        RECT 2.830000 320.380000 4.030000 320.860000 ;
        RECT 7.060000 320.380000 8.260000 320.860000 ;
        RECT 7.060000 331.260000 8.260000 331.740000 ;
        RECT 2.830000 331.260000 4.030000 331.740000 ;
        RECT 2.830000 325.820000 4.030000 326.300000 ;
        RECT 7.060000 325.820000 8.260000 326.300000 ;
        RECT 2.830000 336.700000 4.030000 337.180000 ;
        RECT 7.060000 336.700000 8.260000 337.180000 ;
        RECT 2.830000 342.140000 4.030000 342.620000 ;
        RECT 7.060000 342.140000 8.260000 342.620000 ;
        RECT 2.830000 347.580000 4.030000 348.060000 ;
        RECT 7.060000 347.580000 8.260000 348.060000 ;
        RECT 52.060000 320.380000 53.260000 320.860000 ;
        RECT 52.060000 304.060000 53.260000 304.540000 ;
        RECT 52.060000 309.500000 53.260000 309.980000 ;
        RECT 52.060000 314.940000 53.260000 315.420000 ;
        RECT 97.060000 304.060000 98.260000 304.540000 ;
        RECT 97.060000 309.500000 98.260000 309.980000 ;
        RECT 97.060000 314.940000 98.260000 315.420000 ;
        RECT 97.060000 320.380000 98.260000 320.860000 ;
        RECT 52.060000 325.820000 53.260000 326.300000 ;
        RECT 52.060000 331.260000 53.260000 331.740000 ;
        RECT 52.060000 336.700000 53.260000 337.180000 ;
        RECT 52.060000 342.140000 53.260000 342.620000 ;
        RECT 52.060000 347.580000 53.260000 348.060000 ;
        RECT 97.060000 325.820000 98.260000 326.300000 ;
        RECT 97.060000 331.260000 98.260000 331.740000 ;
        RECT 97.060000 336.700000 98.260000 337.180000 ;
        RECT 97.060000 342.140000 98.260000 342.620000 ;
        RECT 97.060000 347.580000 98.260000 348.060000 ;
        RECT 2.830000 353.020000 4.030000 353.500000 ;
        RECT 7.060000 353.020000 8.260000 353.500000 ;
        RECT 2.830000 358.460000 4.030000 358.940000 ;
        RECT 7.060000 358.460000 8.260000 358.940000 ;
        RECT 2.830000 363.900000 4.030000 364.380000 ;
        RECT 7.060000 363.900000 8.260000 364.380000 ;
        RECT 2.830000 369.340000 4.030000 369.820000 ;
        RECT 2.830000 374.780000 4.030000 375.260000 ;
        RECT 7.060000 369.340000 8.260000 369.820000 ;
        RECT 7.060000 374.780000 8.260000 375.260000 ;
        RECT 2.830000 380.220000 4.030000 380.700000 ;
        RECT 7.060000 380.220000 8.260000 380.700000 ;
        RECT 7.060000 385.660000 8.260000 386.140000 ;
        RECT 2.830000 385.660000 4.030000 386.140000 ;
        RECT 2.830000 391.100000 4.030000 391.580000 ;
        RECT 7.060000 391.100000 8.260000 391.580000 ;
        RECT 52.060000 369.340000 53.260000 369.820000 ;
        RECT 52.060000 353.020000 53.260000 353.500000 ;
        RECT 52.060000 358.460000 53.260000 358.940000 ;
        RECT 52.060000 363.900000 53.260000 364.380000 ;
        RECT 52.060000 374.780000 53.260000 375.260000 ;
        RECT 97.060000 374.780000 98.260000 375.260000 ;
        RECT 97.060000 369.340000 98.260000 369.820000 ;
        RECT 97.060000 353.020000 98.260000 353.500000 ;
        RECT 97.060000 358.460000 98.260000 358.940000 ;
        RECT 97.060000 363.900000 98.260000 364.380000 ;
        RECT 52.060000 380.220000 53.260000 380.700000 ;
        RECT 52.060000 385.660000 53.260000 386.140000 ;
        RECT 52.060000 391.100000 53.260000 391.580000 ;
        RECT 97.060000 380.220000 98.260000 380.700000 ;
        RECT 97.060000 385.660000 98.260000 386.140000 ;
        RECT 97.060000 391.100000 98.260000 391.580000 ;
        RECT 142.060000 222.460000 143.260000 222.940000 ;
        RECT 142.060000 200.700000 143.260000 201.180000 ;
        RECT 142.060000 206.140000 143.260000 206.620000 ;
        RECT 142.060000 211.580000 143.260000 212.060000 ;
        RECT 142.060000 217.020000 143.260000 217.500000 ;
        RECT 142.060000 227.900000 143.260000 228.380000 ;
        RECT 142.060000 233.340000 143.260000 233.820000 ;
        RECT 142.060000 238.780000 143.260000 239.260000 ;
        RECT 142.060000 244.220000 143.260000 244.700000 ;
        RECT 142.060000 249.660000 143.260000 250.140000 ;
        RECT 187.060000 200.700000 188.260000 201.180000 ;
        RECT 187.060000 206.140000 188.260000 206.620000 ;
        RECT 187.060000 211.580000 188.260000 212.060000 ;
        RECT 196.070000 211.580000 197.270000 212.060000 ;
        RECT 196.070000 206.140000 197.270000 206.620000 ;
        RECT 196.070000 200.700000 197.270000 201.180000 ;
        RECT 196.070000 217.020000 197.270000 217.500000 ;
        RECT 196.070000 222.460000 197.270000 222.940000 ;
        RECT 187.060000 222.460000 188.260000 222.940000 ;
        RECT 187.060000 217.020000 188.260000 217.500000 ;
        RECT 196.070000 227.900000 197.270000 228.380000 ;
        RECT 196.070000 233.340000 197.270000 233.820000 ;
        RECT 187.060000 227.900000 188.260000 228.380000 ;
        RECT 187.060000 233.340000 188.260000 233.820000 ;
        RECT 187.060000 238.780000 188.260000 239.260000 ;
        RECT 187.060000 244.220000 188.260000 244.700000 ;
        RECT 187.060000 249.660000 188.260000 250.140000 ;
        RECT 196.070000 249.660000 197.270000 250.140000 ;
        RECT 196.070000 244.220000 197.270000 244.700000 ;
        RECT 196.070000 238.780000 197.270000 239.260000 ;
        RECT 142.060000 271.420000 143.260000 271.900000 ;
        RECT 142.060000 265.980000 143.260000 266.460000 ;
        RECT 142.060000 260.540000 143.260000 261.020000 ;
        RECT 142.060000 255.100000 143.260000 255.580000 ;
        RECT 142.060000 276.860000 143.260000 277.340000 ;
        RECT 142.060000 282.300000 143.260000 282.780000 ;
        RECT 142.060000 287.740000 143.260000 288.220000 ;
        RECT 142.060000 293.180000 143.260000 293.660000 ;
        RECT 142.060000 298.620000 143.260000 299.100000 ;
        RECT 196.070000 255.100000 197.270000 255.580000 ;
        RECT 196.070000 260.540000 197.270000 261.020000 ;
        RECT 187.060000 260.540000 188.260000 261.020000 ;
        RECT 187.060000 255.100000 188.260000 255.580000 ;
        RECT 187.060000 271.420000 188.260000 271.900000 ;
        RECT 187.060000 265.980000 188.260000 266.460000 ;
        RECT 196.070000 271.420000 197.270000 271.900000 ;
        RECT 196.070000 265.980000 197.270000 266.460000 ;
        RECT 196.070000 287.740000 197.270000 288.220000 ;
        RECT 187.060000 287.740000 188.260000 288.220000 ;
        RECT 196.070000 276.860000 197.270000 277.340000 ;
        RECT 196.070000 282.300000 197.270000 282.780000 ;
        RECT 187.060000 276.860000 188.260000 277.340000 ;
        RECT 187.060000 282.300000 188.260000 282.780000 ;
        RECT 196.070000 293.180000 197.270000 293.660000 ;
        RECT 196.070000 298.620000 197.270000 299.100000 ;
        RECT 187.060000 293.180000 188.260000 293.660000 ;
        RECT 187.060000 298.620000 188.260000 299.100000 ;
        RECT 142.060000 320.380000 143.260000 320.860000 ;
        RECT 142.060000 314.940000 143.260000 315.420000 ;
        RECT 142.060000 309.500000 143.260000 309.980000 ;
        RECT 142.060000 304.060000 143.260000 304.540000 ;
        RECT 142.060000 325.820000 143.260000 326.300000 ;
        RECT 142.060000 331.260000 143.260000 331.740000 ;
        RECT 142.060000 336.700000 143.260000 337.180000 ;
        RECT 142.060000 342.140000 143.260000 342.620000 ;
        RECT 142.060000 347.580000 143.260000 348.060000 ;
        RECT 187.060000 309.500000 188.260000 309.980000 ;
        RECT 187.060000 304.060000 188.260000 304.540000 ;
        RECT 196.070000 309.500000 197.270000 309.980000 ;
        RECT 196.070000 304.060000 197.270000 304.540000 ;
        RECT 196.070000 314.940000 197.270000 315.420000 ;
        RECT 196.070000 320.380000 197.270000 320.860000 ;
        RECT 187.060000 320.380000 188.260000 320.860000 ;
        RECT 187.060000 314.940000 188.260000 315.420000 ;
        RECT 187.060000 325.820000 188.260000 326.300000 ;
        RECT 187.060000 331.260000 188.260000 331.740000 ;
        RECT 187.060000 336.700000 188.260000 337.180000 ;
        RECT 196.070000 336.700000 197.270000 337.180000 ;
        RECT 196.070000 331.260000 197.270000 331.740000 ;
        RECT 196.070000 325.820000 197.270000 326.300000 ;
        RECT 196.070000 342.140000 197.270000 342.620000 ;
        RECT 196.070000 347.580000 197.270000 348.060000 ;
        RECT 187.060000 342.140000 188.260000 342.620000 ;
        RECT 187.060000 347.580000 188.260000 348.060000 ;
        RECT 142.060000 369.340000 143.260000 369.820000 ;
        RECT 142.060000 363.900000 143.260000 364.380000 ;
        RECT 142.060000 358.460000 143.260000 358.940000 ;
        RECT 142.060000 353.020000 143.260000 353.500000 ;
        RECT 142.060000 374.780000 143.260000 375.260000 ;
        RECT 142.060000 380.220000 143.260000 380.700000 ;
        RECT 142.060000 385.660000 143.260000 386.140000 ;
        RECT 142.060000 391.100000 143.260000 391.580000 ;
        RECT 196.070000 353.020000 197.270000 353.500000 ;
        RECT 196.070000 358.460000 197.270000 358.940000 ;
        RECT 187.060000 358.460000 188.260000 358.940000 ;
        RECT 187.060000 353.020000 188.260000 353.500000 ;
        RECT 187.060000 369.340000 188.260000 369.820000 ;
        RECT 187.060000 363.900000 188.260000 364.380000 ;
        RECT 187.060000 374.780000 188.260000 375.260000 ;
        RECT 196.070000 374.780000 197.270000 375.260000 ;
        RECT 196.070000 369.340000 197.270000 369.820000 ;
        RECT 196.070000 363.900000 197.270000 364.380000 ;
        RECT 196.070000 380.220000 197.270000 380.700000 ;
        RECT 187.060000 380.220000 188.260000 380.700000 ;
        RECT 187.060000 385.660000 188.260000 386.140000 ;
        RECT 196.070000 385.660000 197.270000 386.140000 ;
        RECT 196.070000 391.100000 197.270000 391.580000 ;
        RECT 187.060000 391.100000 188.260000 391.580000 ;
      LAYER met4 ;
        RECT 187.060000 2.850000 188.260000 396.990000 ;
        RECT 142.060000 2.850000 143.260000 396.990000 ;
        RECT 97.060000 2.850000 98.260000 396.990000 ;
        RECT 52.060000 2.850000 53.260000 396.990000 ;
        RECT 7.060000 2.850000 8.260000 396.990000 ;
        RECT 196.070000 0.000000 197.270000 400.520000 ;
        RECT 2.830000 0.000000 4.030000 400.520000 ;
    END
# end of P/G power stripe data as pin

  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 198.900000 397.590000 200.100000 398.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000000 397.590000 1.200000 398.790000 ;
    END
    PORT
      LAYER met3 ;
        RECT 198.900000 1.050000 200.100000 2.250000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000000 1.050000 1.200000 2.250000 ;
    END
    PORT
      LAYER met4 ;
        RECT 197.870000 399.320000 199.070000 400.520000 ;
    END
    PORT
      LAYER met4 ;
        RECT 197.870000 0.000000 199.070000 1.200000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1.030000 399.320000 2.230000 400.520000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1.030000 0.000000 2.230000 1.200000 ;
    END

# P/G power stripe data as pin
    PORT
      LAYER met3 ;
        RECT 0.000000 1.050000 200.100000 2.250000 ;
        RECT 0.000000 397.590000 200.100000 398.790000 ;
        RECT 4.895000 100.060000 6.260000 100.540000 ;
        RECT 1.030000 100.060000 2.230000 100.540000 ;
        RECT 50.060000 100.060000 51.260000 100.540000 ;
        RECT 95.060000 100.060000 96.260000 100.540000 ;
        RECT 4.895000 7.580000 6.260000 8.060000 ;
        RECT 1.030000 7.580000 2.230000 8.060000 ;
        RECT 4.895000 18.460000 6.260000 18.940000 ;
        RECT 1.030000 18.460000 2.230000 18.940000 ;
        RECT 4.895000 13.020000 6.260000 13.500000 ;
        RECT 1.030000 13.020000 2.230000 13.500000 ;
        RECT 4.895000 23.900000 6.260000 24.380000 ;
        RECT 1.030000 23.900000 2.230000 24.380000 ;
        RECT 4.895000 29.340000 6.260000 29.820000 ;
        RECT 1.030000 29.340000 2.230000 29.820000 ;
        RECT 4.895000 34.780000 6.260000 35.260000 ;
        RECT 1.030000 34.780000 2.230000 35.260000 ;
        RECT 4.895000 40.220000 6.260000 40.700000 ;
        RECT 1.030000 40.220000 2.230000 40.700000 ;
        RECT 4.895000 45.660000 6.260000 46.140000 ;
        RECT 1.030000 45.660000 2.230000 46.140000 ;
        RECT 50.060000 23.900000 51.260000 24.380000 ;
        RECT 50.060000 18.460000 51.260000 18.940000 ;
        RECT 50.060000 13.020000 51.260000 13.500000 ;
        RECT 50.060000 7.580000 51.260000 8.060000 ;
        RECT 95.060000 23.900000 96.260000 24.380000 ;
        RECT 95.060000 18.460000 96.260000 18.940000 ;
        RECT 95.060000 13.020000 96.260000 13.500000 ;
        RECT 95.060000 7.580000 96.260000 8.060000 ;
        RECT 50.060000 45.660000 51.260000 46.140000 ;
        RECT 50.060000 40.220000 51.260000 40.700000 ;
        RECT 50.060000 34.780000 51.260000 35.260000 ;
        RECT 50.060000 29.340000 51.260000 29.820000 ;
        RECT 95.060000 45.660000 96.260000 46.140000 ;
        RECT 95.060000 40.220000 96.260000 40.700000 ;
        RECT 95.060000 34.780000 96.260000 35.260000 ;
        RECT 95.060000 29.340000 96.260000 29.820000 ;
        RECT 4.895000 51.100000 6.260000 51.580000 ;
        RECT 1.030000 51.100000 2.230000 51.580000 ;
        RECT 4.895000 61.980000 6.260000 62.460000 ;
        RECT 1.030000 61.980000 2.230000 62.460000 ;
        RECT 4.895000 56.540000 6.260000 57.020000 ;
        RECT 1.030000 56.540000 2.230000 57.020000 ;
        RECT 4.895000 67.420000 6.260000 67.900000 ;
        RECT 1.030000 67.420000 2.230000 67.900000 ;
        RECT 4.895000 72.860000 6.260000 73.340000 ;
        RECT 1.030000 72.860000 2.230000 73.340000 ;
        RECT 4.895000 78.300000 6.260000 78.780000 ;
        RECT 1.030000 78.300000 2.230000 78.780000 ;
        RECT 4.895000 83.740000 6.260000 84.220000 ;
        RECT 1.030000 83.740000 2.230000 84.220000 ;
        RECT 4.895000 89.180000 6.260000 89.660000 ;
        RECT 1.030000 89.180000 2.230000 89.660000 ;
        RECT 4.895000 94.620000 6.260000 95.100000 ;
        RECT 1.030000 94.620000 2.230000 95.100000 ;
        RECT 50.060000 72.860000 51.260000 73.340000 ;
        RECT 50.060000 67.420000 51.260000 67.900000 ;
        RECT 50.060000 61.980000 51.260000 62.460000 ;
        RECT 50.060000 56.540000 51.260000 57.020000 ;
        RECT 50.060000 51.100000 51.260000 51.580000 ;
        RECT 95.060000 72.860000 96.260000 73.340000 ;
        RECT 95.060000 67.420000 96.260000 67.900000 ;
        RECT 95.060000 61.980000 96.260000 62.460000 ;
        RECT 95.060000 56.540000 96.260000 57.020000 ;
        RECT 95.060000 51.100000 96.260000 51.580000 ;
        RECT 50.060000 94.620000 51.260000 95.100000 ;
        RECT 50.060000 89.180000 51.260000 89.660000 ;
        RECT 50.060000 83.740000 51.260000 84.220000 ;
        RECT 50.060000 78.300000 51.260000 78.780000 ;
        RECT 95.060000 94.620000 96.260000 95.100000 ;
        RECT 95.060000 89.180000 96.260000 89.660000 ;
        RECT 95.060000 83.740000 96.260000 84.220000 ;
        RECT 95.060000 78.300000 96.260000 78.780000 ;
        RECT 4.895000 105.500000 6.260000 105.980000 ;
        RECT 1.030000 105.500000 2.230000 105.980000 ;
        RECT 4.895000 110.940000 6.260000 111.420000 ;
        RECT 1.030000 110.940000 2.230000 111.420000 ;
        RECT 4.895000 116.380000 6.260000 116.860000 ;
        RECT 1.030000 116.380000 2.230000 116.860000 ;
        RECT 4.895000 121.820000 6.260000 122.300000 ;
        RECT 1.030000 121.820000 2.230000 122.300000 ;
        RECT 4.895000 127.260000 6.260000 127.740000 ;
        RECT 1.030000 127.260000 2.230000 127.740000 ;
        RECT 4.895000 132.700000 6.260000 133.180000 ;
        RECT 1.030000 132.700000 2.230000 133.180000 ;
        RECT 4.895000 143.580000 6.260000 144.060000 ;
        RECT 1.030000 143.580000 2.230000 144.060000 ;
        RECT 4.895000 138.140000 6.260000 138.620000 ;
        RECT 1.030000 138.140000 2.230000 138.620000 ;
        RECT 4.895000 149.020000 6.260000 149.500000 ;
        RECT 1.030000 149.020000 2.230000 149.500000 ;
        RECT 50.060000 121.820000 51.260000 122.300000 ;
        RECT 50.060000 116.380000 51.260000 116.860000 ;
        RECT 50.060000 110.940000 51.260000 111.420000 ;
        RECT 50.060000 105.500000 51.260000 105.980000 ;
        RECT 95.060000 121.820000 96.260000 122.300000 ;
        RECT 95.060000 116.380000 96.260000 116.860000 ;
        RECT 95.060000 110.940000 96.260000 111.420000 ;
        RECT 95.060000 105.500000 96.260000 105.980000 ;
        RECT 50.060000 149.020000 51.260000 149.500000 ;
        RECT 50.060000 143.580000 51.260000 144.060000 ;
        RECT 50.060000 138.140000 51.260000 138.620000 ;
        RECT 50.060000 132.700000 51.260000 133.180000 ;
        RECT 50.060000 127.260000 51.260000 127.740000 ;
        RECT 95.060000 149.020000 96.260000 149.500000 ;
        RECT 95.060000 143.580000 96.260000 144.060000 ;
        RECT 95.060000 138.140000 96.260000 138.620000 ;
        RECT 95.060000 132.700000 96.260000 133.180000 ;
        RECT 95.060000 127.260000 96.260000 127.740000 ;
        RECT 4.895000 154.460000 6.260000 154.940000 ;
        RECT 1.030000 154.460000 2.230000 154.940000 ;
        RECT 4.895000 159.900000 6.260000 160.380000 ;
        RECT 1.030000 159.900000 2.230000 160.380000 ;
        RECT 4.895000 165.340000 6.260000 165.820000 ;
        RECT 1.030000 165.340000 2.230000 165.820000 ;
        RECT 4.895000 170.780000 6.260000 171.260000 ;
        RECT 1.030000 170.780000 2.230000 171.260000 ;
        RECT 4.895000 176.220000 6.260000 176.700000 ;
        RECT 1.030000 176.220000 2.230000 176.700000 ;
        RECT 4.895000 187.100000 6.260000 187.580000 ;
        RECT 1.030000 187.100000 2.230000 187.580000 ;
        RECT 4.895000 181.660000 6.260000 182.140000 ;
        RECT 1.030000 181.660000 2.230000 182.140000 ;
        RECT 4.895000 192.540000 6.260000 193.020000 ;
        RECT 1.030000 192.540000 2.230000 193.020000 ;
        RECT 4.895000 197.980000 6.260000 198.460000 ;
        RECT 1.030000 197.980000 2.230000 198.460000 ;
        RECT 50.060000 170.780000 51.260000 171.260000 ;
        RECT 50.060000 165.340000 51.260000 165.820000 ;
        RECT 50.060000 159.900000 51.260000 160.380000 ;
        RECT 50.060000 154.460000 51.260000 154.940000 ;
        RECT 95.060000 170.780000 96.260000 171.260000 ;
        RECT 95.060000 165.340000 96.260000 165.820000 ;
        RECT 95.060000 159.900000 96.260000 160.380000 ;
        RECT 95.060000 154.460000 96.260000 154.940000 ;
        RECT 50.060000 197.980000 51.260000 198.460000 ;
        RECT 50.060000 192.540000 51.260000 193.020000 ;
        RECT 50.060000 187.100000 51.260000 187.580000 ;
        RECT 50.060000 181.660000 51.260000 182.140000 ;
        RECT 50.060000 176.220000 51.260000 176.700000 ;
        RECT 95.060000 197.980000 96.260000 198.460000 ;
        RECT 95.060000 192.540000 96.260000 193.020000 ;
        RECT 95.060000 187.100000 96.260000 187.580000 ;
        RECT 95.060000 181.660000 96.260000 182.140000 ;
        RECT 95.060000 176.220000 96.260000 176.700000 ;
        RECT 197.870000 100.060000 199.070000 100.540000 ;
        RECT 140.060000 100.060000 141.260000 100.540000 ;
        RECT 185.060000 100.060000 186.260000 100.540000 ;
        RECT 140.060000 23.900000 141.260000 24.380000 ;
        RECT 140.060000 18.460000 141.260000 18.940000 ;
        RECT 140.060000 13.020000 141.260000 13.500000 ;
        RECT 140.060000 7.580000 141.260000 8.060000 ;
        RECT 140.060000 45.660000 141.260000 46.140000 ;
        RECT 140.060000 40.220000 141.260000 40.700000 ;
        RECT 140.060000 34.780000 141.260000 35.260000 ;
        RECT 140.060000 29.340000 141.260000 29.820000 ;
        RECT 197.870000 7.580000 199.070000 8.060000 ;
        RECT 185.060000 7.580000 186.260000 8.060000 ;
        RECT 185.060000 13.020000 186.260000 13.500000 ;
        RECT 185.060000 18.460000 186.260000 18.940000 ;
        RECT 185.060000 23.900000 186.260000 24.380000 ;
        RECT 197.870000 23.900000 199.070000 24.380000 ;
        RECT 197.870000 13.020000 199.070000 13.500000 ;
        RECT 197.870000 18.460000 199.070000 18.940000 ;
        RECT 197.870000 34.780000 199.070000 35.260000 ;
        RECT 197.870000 29.340000 199.070000 29.820000 ;
        RECT 185.060000 34.780000 186.260000 35.260000 ;
        RECT 185.060000 29.340000 186.260000 29.820000 ;
        RECT 197.870000 45.660000 199.070000 46.140000 ;
        RECT 197.870000 40.220000 199.070000 40.700000 ;
        RECT 185.060000 45.660000 186.260000 46.140000 ;
        RECT 185.060000 40.220000 186.260000 40.700000 ;
        RECT 140.060000 72.860000 141.260000 73.340000 ;
        RECT 140.060000 67.420000 141.260000 67.900000 ;
        RECT 140.060000 61.980000 141.260000 62.460000 ;
        RECT 140.060000 56.540000 141.260000 57.020000 ;
        RECT 140.060000 51.100000 141.260000 51.580000 ;
        RECT 140.060000 94.620000 141.260000 95.100000 ;
        RECT 140.060000 89.180000 141.260000 89.660000 ;
        RECT 140.060000 83.740000 141.260000 84.220000 ;
        RECT 140.060000 78.300000 141.260000 78.780000 ;
        RECT 185.060000 51.100000 186.260000 51.580000 ;
        RECT 185.060000 56.540000 186.260000 57.020000 ;
        RECT 185.060000 61.980000 186.260000 62.460000 ;
        RECT 197.870000 61.980000 199.070000 62.460000 ;
        RECT 197.870000 51.100000 199.070000 51.580000 ;
        RECT 197.870000 56.540000 199.070000 57.020000 ;
        RECT 197.870000 72.860000 199.070000 73.340000 ;
        RECT 197.870000 67.420000 199.070000 67.900000 ;
        RECT 185.060000 72.860000 186.260000 73.340000 ;
        RECT 185.060000 67.420000 186.260000 67.900000 ;
        RECT 185.060000 78.300000 186.260000 78.780000 ;
        RECT 185.060000 83.740000 186.260000 84.220000 ;
        RECT 197.870000 83.740000 199.070000 84.220000 ;
        RECT 197.870000 78.300000 199.070000 78.780000 ;
        RECT 197.870000 94.620000 199.070000 95.100000 ;
        RECT 197.870000 89.180000 199.070000 89.660000 ;
        RECT 185.060000 94.620000 186.260000 95.100000 ;
        RECT 185.060000 89.180000 186.260000 89.660000 ;
        RECT 140.060000 121.820000 141.260000 122.300000 ;
        RECT 140.060000 116.380000 141.260000 116.860000 ;
        RECT 140.060000 110.940000 141.260000 111.420000 ;
        RECT 140.060000 105.500000 141.260000 105.980000 ;
        RECT 140.060000 149.020000 141.260000 149.500000 ;
        RECT 140.060000 143.580000 141.260000 144.060000 ;
        RECT 140.060000 138.140000 141.260000 138.620000 ;
        RECT 140.060000 132.700000 141.260000 133.180000 ;
        RECT 140.060000 127.260000 141.260000 127.740000 ;
        RECT 197.870000 110.940000 199.070000 111.420000 ;
        RECT 197.870000 105.500000 199.070000 105.980000 ;
        RECT 185.060000 110.940000 186.260000 111.420000 ;
        RECT 185.060000 105.500000 186.260000 105.980000 ;
        RECT 185.060000 116.380000 186.260000 116.860000 ;
        RECT 185.060000 121.820000 186.260000 122.300000 ;
        RECT 197.870000 121.820000 199.070000 122.300000 ;
        RECT 197.870000 116.380000 199.070000 116.860000 ;
        RECT 197.870000 132.700000 199.070000 133.180000 ;
        RECT 197.870000 127.260000 199.070000 127.740000 ;
        RECT 185.060000 132.700000 186.260000 133.180000 ;
        RECT 185.060000 127.260000 186.260000 127.740000 ;
        RECT 185.060000 138.140000 186.260000 138.620000 ;
        RECT 185.060000 143.580000 186.260000 144.060000 ;
        RECT 185.060000 149.020000 186.260000 149.500000 ;
        RECT 197.870000 149.020000 199.070000 149.500000 ;
        RECT 197.870000 138.140000 199.070000 138.620000 ;
        RECT 197.870000 143.580000 199.070000 144.060000 ;
        RECT 140.060000 170.780000 141.260000 171.260000 ;
        RECT 140.060000 165.340000 141.260000 165.820000 ;
        RECT 140.060000 159.900000 141.260000 160.380000 ;
        RECT 140.060000 154.460000 141.260000 154.940000 ;
        RECT 140.060000 197.980000 141.260000 198.460000 ;
        RECT 140.060000 192.540000 141.260000 193.020000 ;
        RECT 140.060000 187.100000 141.260000 187.580000 ;
        RECT 140.060000 181.660000 141.260000 182.140000 ;
        RECT 140.060000 176.220000 141.260000 176.700000 ;
        RECT 197.870000 159.900000 199.070000 160.380000 ;
        RECT 197.870000 154.460000 199.070000 154.940000 ;
        RECT 185.060000 159.900000 186.260000 160.380000 ;
        RECT 185.060000 154.460000 186.260000 154.940000 ;
        RECT 197.870000 170.780000 199.070000 171.260000 ;
        RECT 197.870000 165.340000 199.070000 165.820000 ;
        RECT 185.060000 170.780000 186.260000 171.260000 ;
        RECT 185.060000 165.340000 186.260000 165.820000 ;
        RECT 185.060000 176.220000 186.260000 176.700000 ;
        RECT 185.060000 181.660000 186.260000 182.140000 ;
        RECT 185.060000 187.100000 186.260000 187.580000 ;
        RECT 197.870000 187.100000 199.070000 187.580000 ;
        RECT 197.870000 176.220000 199.070000 176.700000 ;
        RECT 197.870000 181.660000 199.070000 182.140000 ;
        RECT 197.870000 197.980000 199.070000 198.460000 ;
        RECT 197.870000 192.540000 199.070000 193.020000 ;
        RECT 185.060000 197.980000 186.260000 198.460000 ;
        RECT 185.060000 192.540000 186.260000 193.020000 ;
        RECT 4.895000 225.180000 6.260000 225.660000 ;
        RECT 1.030000 225.180000 2.230000 225.660000 ;
        RECT 4.895000 203.420000 6.260000 203.900000 ;
        RECT 1.030000 203.420000 2.230000 203.900000 ;
        RECT 4.895000 208.860000 6.260000 209.340000 ;
        RECT 1.030000 208.860000 2.230000 209.340000 ;
        RECT 4.895000 214.300000 6.260000 214.780000 ;
        RECT 1.030000 214.300000 2.230000 214.780000 ;
        RECT 4.895000 219.740000 6.260000 220.220000 ;
        RECT 1.030000 219.740000 2.230000 220.220000 ;
        RECT 4.895000 230.620000 6.260000 231.100000 ;
        RECT 1.030000 230.620000 2.230000 231.100000 ;
        RECT 4.895000 236.060000 6.260000 236.540000 ;
        RECT 1.030000 236.060000 2.230000 236.540000 ;
        RECT 4.895000 241.500000 6.260000 241.980000 ;
        RECT 1.030000 241.500000 2.230000 241.980000 ;
        RECT 4.895000 246.940000 6.260000 247.420000 ;
        RECT 1.030000 246.940000 2.230000 247.420000 ;
        RECT 50.060000 225.180000 51.260000 225.660000 ;
        RECT 95.060000 225.180000 96.260000 225.660000 ;
        RECT 50.060000 219.740000 51.260000 220.220000 ;
        RECT 50.060000 214.300000 51.260000 214.780000 ;
        RECT 50.060000 208.860000 51.260000 209.340000 ;
        RECT 50.060000 203.420000 51.260000 203.900000 ;
        RECT 95.060000 219.740000 96.260000 220.220000 ;
        RECT 95.060000 214.300000 96.260000 214.780000 ;
        RECT 95.060000 208.860000 96.260000 209.340000 ;
        RECT 95.060000 203.420000 96.260000 203.900000 ;
        RECT 50.060000 246.940000 51.260000 247.420000 ;
        RECT 50.060000 241.500000 51.260000 241.980000 ;
        RECT 50.060000 236.060000 51.260000 236.540000 ;
        RECT 50.060000 230.620000 51.260000 231.100000 ;
        RECT 95.060000 246.940000 96.260000 247.420000 ;
        RECT 95.060000 241.500000 96.260000 241.980000 ;
        RECT 95.060000 236.060000 96.260000 236.540000 ;
        RECT 95.060000 230.620000 96.260000 231.100000 ;
        RECT 4.895000 252.380000 6.260000 252.860000 ;
        RECT 1.030000 252.380000 2.230000 252.860000 ;
        RECT 4.895000 257.820000 6.260000 258.300000 ;
        RECT 1.030000 257.820000 2.230000 258.300000 ;
        RECT 4.895000 268.700000 6.260000 269.180000 ;
        RECT 1.030000 268.700000 2.230000 269.180000 ;
        RECT 4.895000 263.260000 6.260000 263.740000 ;
        RECT 1.030000 263.260000 2.230000 263.740000 ;
        RECT 4.895000 274.140000 6.260000 274.620000 ;
        RECT 1.030000 274.140000 2.230000 274.620000 ;
        RECT 4.895000 279.580000 6.260000 280.060000 ;
        RECT 1.030000 279.580000 2.230000 280.060000 ;
        RECT 4.895000 285.020000 6.260000 285.500000 ;
        RECT 1.030000 285.020000 2.230000 285.500000 ;
        RECT 4.895000 290.460000 6.260000 290.940000 ;
        RECT 1.030000 290.460000 2.230000 290.940000 ;
        RECT 4.895000 295.900000 6.260000 296.380000 ;
        RECT 1.030000 295.900000 2.230000 296.380000 ;
        RECT 50.060000 274.140000 51.260000 274.620000 ;
        RECT 50.060000 268.700000 51.260000 269.180000 ;
        RECT 50.060000 263.260000 51.260000 263.740000 ;
        RECT 50.060000 257.820000 51.260000 258.300000 ;
        RECT 50.060000 252.380000 51.260000 252.860000 ;
        RECT 95.060000 274.140000 96.260000 274.620000 ;
        RECT 95.060000 268.700000 96.260000 269.180000 ;
        RECT 95.060000 263.260000 96.260000 263.740000 ;
        RECT 95.060000 257.820000 96.260000 258.300000 ;
        RECT 95.060000 252.380000 96.260000 252.860000 ;
        RECT 50.060000 295.900000 51.260000 296.380000 ;
        RECT 50.060000 290.460000 51.260000 290.940000 ;
        RECT 50.060000 285.020000 51.260000 285.500000 ;
        RECT 50.060000 279.580000 51.260000 280.060000 ;
        RECT 95.060000 295.900000 96.260000 296.380000 ;
        RECT 95.060000 290.460000 96.260000 290.940000 ;
        RECT 95.060000 285.020000 96.260000 285.500000 ;
        RECT 95.060000 279.580000 96.260000 280.060000 ;
        RECT 4.895000 350.300000 6.260000 350.780000 ;
        RECT 1.030000 350.300000 2.230000 350.780000 ;
        RECT 50.060000 350.300000 51.260000 350.780000 ;
        RECT 95.060000 350.300000 96.260000 350.780000 ;
        RECT 4.895000 301.340000 6.260000 301.820000 ;
        RECT 1.030000 301.340000 2.230000 301.820000 ;
        RECT 4.895000 312.220000 6.260000 312.700000 ;
        RECT 1.030000 312.220000 2.230000 312.700000 ;
        RECT 4.895000 306.780000 6.260000 307.260000 ;
        RECT 1.030000 306.780000 2.230000 307.260000 ;
        RECT 4.895000 317.660000 6.260000 318.140000 ;
        RECT 1.030000 317.660000 2.230000 318.140000 ;
        RECT 4.895000 323.100000 6.260000 323.580000 ;
        RECT 1.030000 323.100000 2.230000 323.580000 ;
        RECT 4.895000 328.540000 6.260000 329.020000 ;
        RECT 1.030000 328.540000 2.230000 329.020000 ;
        RECT 4.895000 333.980000 6.260000 334.460000 ;
        RECT 1.030000 333.980000 2.230000 334.460000 ;
        RECT 4.895000 339.420000 6.260000 339.900000 ;
        RECT 1.030000 339.420000 2.230000 339.900000 ;
        RECT 4.895000 344.860000 6.260000 345.340000 ;
        RECT 1.030000 344.860000 2.230000 345.340000 ;
        RECT 50.060000 323.100000 51.260000 323.580000 ;
        RECT 50.060000 317.660000 51.260000 318.140000 ;
        RECT 50.060000 312.220000 51.260000 312.700000 ;
        RECT 50.060000 306.780000 51.260000 307.260000 ;
        RECT 50.060000 301.340000 51.260000 301.820000 ;
        RECT 95.060000 323.100000 96.260000 323.580000 ;
        RECT 95.060000 317.660000 96.260000 318.140000 ;
        RECT 95.060000 312.220000 96.260000 312.700000 ;
        RECT 95.060000 306.780000 96.260000 307.260000 ;
        RECT 95.060000 301.340000 96.260000 301.820000 ;
        RECT 50.060000 344.860000 51.260000 345.340000 ;
        RECT 50.060000 339.420000 51.260000 339.900000 ;
        RECT 50.060000 333.980000 51.260000 334.460000 ;
        RECT 50.060000 328.540000 51.260000 329.020000 ;
        RECT 95.060000 344.860000 96.260000 345.340000 ;
        RECT 95.060000 339.420000 96.260000 339.900000 ;
        RECT 95.060000 333.980000 96.260000 334.460000 ;
        RECT 95.060000 328.540000 96.260000 329.020000 ;
        RECT 4.895000 355.740000 6.260000 356.220000 ;
        RECT 1.030000 355.740000 2.230000 356.220000 ;
        RECT 4.895000 361.180000 6.260000 361.660000 ;
        RECT 1.030000 361.180000 2.230000 361.660000 ;
        RECT 4.895000 366.620000 6.260000 367.100000 ;
        RECT 1.030000 366.620000 2.230000 367.100000 ;
        RECT 4.895000 372.060000 6.260000 372.540000 ;
        RECT 1.030000 372.060000 2.230000 372.540000 ;
        RECT 4.895000 377.500000 6.260000 377.980000 ;
        RECT 1.030000 377.500000 2.230000 377.980000 ;
        RECT 4.895000 382.940000 6.260000 383.420000 ;
        RECT 1.030000 382.940000 2.230000 383.420000 ;
        RECT 4.895000 393.820000 6.260000 394.300000 ;
        RECT 1.030000 393.820000 2.230000 394.300000 ;
        RECT 4.895000 388.380000 6.260000 388.860000 ;
        RECT 1.030000 388.380000 2.230000 388.860000 ;
        RECT 50.060000 372.060000 51.260000 372.540000 ;
        RECT 50.060000 366.620000 51.260000 367.100000 ;
        RECT 50.060000 361.180000 51.260000 361.660000 ;
        RECT 50.060000 355.740000 51.260000 356.220000 ;
        RECT 95.060000 372.060000 96.260000 372.540000 ;
        RECT 95.060000 366.620000 96.260000 367.100000 ;
        RECT 95.060000 361.180000 96.260000 361.660000 ;
        RECT 95.060000 355.740000 96.260000 356.220000 ;
        RECT 50.060000 393.820000 51.260000 394.300000 ;
        RECT 50.060000 388.380000 51.260000 388.860000 ;
        RECT 50.060000 382.940000 51.260000 383.420000 ;
        RECT 50.060000 377.500000 51.260000 377.980000 ;
        RECT 95.060000 393.820000 96.260000 394.300000 ;
        RECT 95.060000 388.380000 96.260000 388.860000 ;
        RECT 95.060000 377.500000 96.260000 377.980000 ;
        RECT 95.060000 382.940000 96.260000 383.420000 ;
        RECT 140.060000 225.180000 141.260000 225.660000 ;
        RECT 140.060000 219.740000 141.260000 220.220000 ;
        RECT 140.060000 214.300000 141.260000 214.780000 ;
        RECT 140.060000 208.860000 141.260000 209.340000 ;
        RECT 140.060000 203.420000 141.260000 203.900000 ;
        RECT 140.060000 246.940000 141.260000 247.420000 ;
        RECT 140.060000 241.500000 141.260000 241.980000 ;
        RECT 140.060000 236.060000 141.260000 236.540000 ;
        RECT 140.060000 230.620000 141.260000 231.100000 ;
        RECT 197.870000 225.180000 199.070000 225.660000 ;
        RECT 185.060000 225.180000 186.260000 225.660000 ;
        RECT 185.060000 203.420000 186.260000 203.900000 ;
        RECT 185.060000 208.860000 186.260000 209.340000 ;
        RECT 197.870000 208.860000 199.070000 209.340000 ;
        RECT 197.870000 203.420000 199.070000 203.900000 ;
        RECT 197.870000 219.740000 199.070000 220.220000 ;
        RECT 197.870000 214.300000 199.070000 214.780000 ;
        RECT 185.060000 219.740000 186.260000 220.220000 ;
        RECT 185.060000 214.300000 186.260000 214.780000 ;
        RECT 197.870000 236.060000 199.070000 236.540000 ;
        RECT 197.870000 230.620000 199.070000 231.100000 ;
        RECT 185.060000 236.060000 186.260000 236.540000 ;
        RECT 185.060000 230.620000 186.260000 231.100000 ;
        RECT 185.060000 241.500000 186.260000 241.980000 ;
        RECT 185.060000 246.940000 186.260000 247.420000 ;
        RECT 197.870000 246.940000 199.070000 247.420000 ;
        RECT 197.870000 241.500000 199.070000 241.980000 ;
        RECT 140.060000 274.140000 141.260000 274.620000 ;
        RECT 140.060000 268.700000 141.260000 269.180000 ;
        RECT 140.060000 263.260000 141.260000 263.740000 ;
        RECT 140.060000 257.820000 141.260000 258.300000 ;
        RECT 140.060000 252.380000 141.260000 252.860000 ;
        RECT 140.060000 295.900000 141.260000 296.380000 ;
        RECT 140.060000 290.460000 141.260000 290.940000 ;
        RECT 140.060000 285.020000 141.260000 285.500000 ;
        RECT 140.060000 279.580000 141.260000 280.060000 ;
        RECT 197.870000 257.820000 199.070000 258.300000 ;
        RECT 197.870000 252.380000 199.070000 252.860000 ;
        RECT 185.060000 257.820000 186.260000 258.300000 ;
        RECT 185.060000 252.380000 186.260000 252.860000 ;
        RECT 185.060000 263.260000 186.260000 263.740000 ;
        RECT 185.060000 268.700000 186.260000 269.180000 ;
        RECT 185.060000 274.140000 186.260000 274.620000 ;
        RECT 197.870000 274.140000 199.070000 274.620000 ;
        RECT 197.870000 263.260000 199.070000 263.740000 ;
        RECT 197.870000 268.700000 199.070000 269.180000 ;
        RECT 197.870000 285.020000 199.070000 285.500000 ;
        RECT 197.870000 279.580000 199.070000 280.060000 ;
        RECT 185.060000 285.020000 186.260000 285.500000 ;
        RECT 185.060000 279.580000 186.260000 280.060000 ;
        RECT 197.870000 295.900000 199.070000 296.380000 ;
        RECT 197.870000 290.460000 199.070000 290.940000 ;
        RECT 185.060000 295.900000 186.260000 296.380000 ;
        RECT 185.060000 290.460000 186.260000 290.940000 ;
        RECT 197.870000 350.300000 199.070000 350.780000 ;
        RECT 140.060000 350.300000 141.260000 350.780000 ;
        RECT 185.060000 350.300000 186.260000 350.780000 ;
        RECT 140.060000 323.100000 141.260000 323.580000 ;
        RECT 140.060000 317.660000 141.260000 318.140000 ;
        RECT 140.060000 312.220000 141.260000 312.700000 ;
        RECT 140.060000 306.780000 141.260000 307.260000 ;
        RECT 140.060000 301.340000 141.260000 301.820000 ;
        RECT 140.060000 344.860000 141.260000 345.340000 ;
        RECT 140.060000 339.420000 141.260000 339.900000 ;
        RECT 140.060000 333.980000 141.260000 334.460000 ;
        RECT 140.060000 328.540000 141.260000 329.020000 ;
        RECT 185.060000 301.340000 186.260000 301.820000 ;
        RECT 185.060000 306.780000 186.260000 307.260000 ;
        RECT 185.060000 312.220000 186.260000 312.700000 ;
        RECT 197.870000 312.220000 199.070000 312.700000 ;
        RECT 197.870000 301.340000 199.070000 301.820000 ;
        RECT 197.870000 306.780000 199.070000 307.260000 ;
        RECT 197.870000 323.100000 199.070000 323.580000 ;
        RECT 197.870000 317.660000 199.070000 318.140000 ;
        RECT 185.060000 323.100000 186.260000 323.580000 ;
        RECT 185.060000 317.660000 186.260000 318.140000 ;
        RECT 185.060000 328.540000 186.260000 329.020000 ;
        RECT 185.060000 333.980000 186.260000 334.460000 ;
        RECT 197.870000 333.980000 199.070000 334.460000 ;
        RECT 197.870000 328.540000 199.070000 329.020000 ;
        RECT 197.870000 344.860000 199.070000 345.340000 ;
        RECT 197.870000 339.420000 199.070000 339.900000 ;
        RECT 185.060000 344.860000 186.260000 345.340000 ;
        RECT 185.060000 339.420000 186.260000 339.900000 ;
        RECT 140.060000 372.060000 141.260000 372.540000 ;
        RECT 140.060000 366.620000 141.260000 367.100000 ;
        RECT 140.060000 355.740000 141.260000 356.220000 ;
        RECT 140.060000 361.180000 141.260000 361.660000 ;
        RECT 140.060000 393.820000 141.260000 394.300000 ;
        RECT 140.060000 388.380000 141.260000 388.860000 ;
        RECT 140.060000 382.940000 141.260000 383.420000 ;
        RECT 140.060000 377.500000 141.260000 377.980000 ;
        RECT 197.870000 361.180000 199.070000 361.660000 ;
        RECT 197.870000 355.740000 199.070000 356.220000 ;
        RECT 185.060000 361.180000 186.260000 361.660000 ;
        RECT 185.060000 355.740000 186.260000 356.220000 ;
        RECT 185.060000 366.620000 186.260000 367.100000 ;
        RECT 185.060000 372.060000 186.260000 372.540000 ;
        RECT 197.870000 372.060000 199.070000 372.540000 ;
        RECT 197.870000 366.620000 199.070000 367.100000 ;
        RECT 197.870000 382.940000 199.070000 383.420000 ;
        RECT 197.870000 377.500000 199.070000 377.980000 ;
        RECT 185.060000 382.940000 186.260000 383.420000 ;
        RECT 185.060000 377.500000 186.260000 377.980000 ;
        RECT 197.870000 393.820000 199.070000 394.300000 ;
        RECT 197.870000 388.380000 199.070000 388.860000 ;
        RECT 185.060000 393.820000 186.260000 394.300000 ;
        RECT 185.060000 388.380000 186.260000 388.860000 ;
      LAYER met4 ;
        RECT 185.060000 1.050000 186.260000 398.790000 ;
        RECT 140.060000 1.050000 141.260000 398.790000 ;
        RECT 95.060000 1.050000 96.260000 398.790000 ;
        RECT 50.060000 1.050000 51.260000 398.790000 ;
        RECT 5.060000 1.050000 6.260000 398.790000 ;
        RECT 197.870000 0.000000 199.070000 400.520000 ;
        RECT 1.030000 0.000000 2.230000 400.520000 ;
        RECT 4.895000 100.060000 6.260000 100.540000 ;
        RECT 4.895000 7.580000 6.260000 8.060000 ;
        RECT 4.895000 18.460000 6.260000 18.940000 ;
        RECT 4.895000 13.020000 6.260000 13.500000 ;
        RECT 4.895000 23.900000 6.260000 24.380000 ;
        RECT 4.895000 29.340000 6.260000 29.820000 ;
        RECT 4.895000 34.780000 6.260000 35.260000 ;
        RECT 4.895000 40.220000 6.260000 40.700000 ;
        RECT 4.895000 45.660000 6.260000 46.140000 ;
        RECT 4.895000 51.100000 6.260000 51.580000 ;
        RECT 4.895000 61.980000 6.260000 62.460000 ;
        RECT 4.895000 56.540000 6.260000 57.020000 ;
        RECT 4.895000 67.420000 6.260000 67.900000 ;
        RECT 4.895000 72.860000 6.260000 73.340000 ;
        RECT 4.895000 78.300000 6.260000 78.780000 ;
        RECT 4.895000 83.740000 6.260000 84.220000 ;
        RECT 4.895000 89.180000 6.260000 89.660000 ;
        RECT 4.895000 94.620000 6.260000 95.100000 ;
        RECT 4.895000 105.500000 6.260000 105.980000 ;
        RECT 4.895000 110.940000 6.260000 111.420000 ;
        RECT 4.895000 116.380000 6.260000 116.860000 ;
        RECT 4.895000 121.820000 6.260000 122.300000 ;
        RECT 4.895000 127.260000 6.260000 127.740000 ;
        RECT 4.895000 132.700000 6.260000 133.180000 ;
        RECT 4.895000 143.580000 6.260000 144.060000 ;
        RECT 4.895000 138.140000 6.260000 138.620000 ;
        RECT 4.895000 149.020000 6.260000 149.500000 ;
        RECT 4.895000 154.460000 6.260000 154.940000 ;
        RECT 4.895000 159.900000 6.260000 160.380000 ;
        RECT 4.895000 165.340000 6.260000 165.820000 ;
        RECT 4.895000 170.780000 6.260000 171.260000 ;
        RECT 4.895000 176.220000 6.260000 176.700000 ;
        RECT 4.895000 187.100000 6.260000 187.580000 ;
        RECT 4.895000 181.660000 6.260000 182.140000 ;
        RECT 4.895000 192.540000 6.260000 193.020000 ;
        RECT 4.895000 197.980000 6.260000 198.460000 ;
        RECT 4.895000 225.180000 6.260000 225.660000 ;
        RECT 4.895000 203.420000 6.260000 203.900000 ;
        RECT 4.895000 208.860000 6.260000 209.340000 ;
        RECT 4.895000 214.300000 6.260000 214.780000 ;
        RECT 4.895000 219.740000 6.260000 220.220000 ;
        RECT 4.895000 230.620000 6.260000 231.100000 ;
        RECT 4.895000 236.060000 6.260000 236.540000 ;
        RECT 4.895000 241.500000 6.260000 241.980000 ;
        RECT 4.895000 246.940000 6.260000 247.420000 ;
        RECT 4.895000 252.380000 6.260000 252.860000 ;
        RECT 4.895000 257.820000 6.260000 258.300000 ;
        RECT 4.895000 268.700000 6.260000 269.180000 ;
        RECT 4.895000 263.260000 6.260000 263.740000 ;
        RECT 4.895000 274.140000 6.260000 274.620000 ;
        RECT 4.895000 279.580000 6.260000 280.060000 ;
        RECT 4.895000 285.020000 6.260000 285.500000 ;
        RECT 4.895000 290.460000 6.260000 290.940000 ;
        RECT 4.895000 295.900000 6.260000 296.380000 ;
        RECT 4.895000 350.300000 6.260000 350.780000 ;
        RECT 4.895000 301.340000 6.260000 301.820000 ;
        RECT 4.895000 312.220000 6.260000 312.700000 ;
        RECT 4.895000 306.780000 6.260000 307.260000 ;
        RECT 4.895000 317.660000 6.260000 318.140000 ;
        RECT 4.895000 323.100000 6.260000 323.580000 ;
        RECT 4.895000 328.540000 6.260000 329.020000 ;
        RECT 4.895000 333.980000 6.260000 334.460000 ;
        RECT 4.895000 339.420000 6.260000 339.900000 ;
        RECT 4.895000 344.860000 6.260000 345.340000 ;
        RECT 4.895000 355.740000 6.260000 356.220000 ;
        RECT 4.895000 361.180000 6.260000 361.660000 ;
        RECT 4.895000 366.620000 6.260000 367.100000 ;
        RECT 4.895000 372.060000 6.260000 372.540000 ;
        RECT 4.895000 377.500000 6.260000 377.980000 ;
        RECT 4.895000 382.940000 6.260000 383.420000 ;
        RECT 4.895000 393.820000 6.260000 394.300000 ;
        RECT 4.895000 388.380000 6.260000 388.860000 ;
    END
# end of P/G power stripe data as pin

  END vssd1
  OBS
    LAYER li1 ;
      RECT 0.000000 0.000000 200.100000 400.520000 ;
    LAYER met1 ;
      RECT 0.000000 0.000000 200.100000 400.520000 ;
    LAYER met2 ;
      RECT 194.680000 399.680000 200.100000 400.520000 ;
      RECT 193.300000 399.680000 194.020000 400.520000 ;
      RECT 191.920000 399.680000 192.640000 400.520000 ;
      RECT 190.540000 399.680000 191.260000 400.520000 ;
      RECT 188.700000 399.680000 189.880000 400.520000 ;
      RECT 187.320000 399.680000 188.040000 400.520000 ;
      RECT 185.940000 399.680000 186.660000 400.520000 ;
      RECT 184.100000 399.680000 185.280000 400.520000 ;
      RECT 182.720000 399.680000 183.440000 400.520000 ;
      RECT 181.340000 399.680000 182.060000 400.520000 ;
      RECT 179.500000 399.680000 180.680000 400.520000 ;
      RECT 178.120000 399.680000 178.840000 400.520000 ;
      RECT 176.740000 399.680000 177.460000 400.520000 ;
      RECT 174.900000 399.680000 176.080000 400.520000 ;
      RECT 173.520000 399.680000 174.240000 400.520000 ;
      RECT 172.140000 399.680000 172.860000 400.520000 ;
      RECT 170.300000 399.680000 171.480000 400.520000 ;
      RECT 168.920000 399.680000 169.640000 400.520000 ;
      RECT 167.540000 399.680000 168.260000 400.520000 ;
      RECT 165.700000 399.680000 166.880000 400.520000 ;
      RECT 164.320000 399.680000 165.040000 400.520000 ;
      RECT 162.940000 399.680000 163.660000 400.520000 ;
      RECT 161.100000 399.680000 162.280000 400.520000 ;
      RECT 159.720000 399.680000 160.440000 400.520000 ;
      RECT 158.340000 399.680000 159.060000 400.520000 ;
      RECT 156.500000 399.680000 157.680000 400.520000 ;
      RECT 155.120000 399.680000 155.840000 400.520000 ;
      RECT 153.740000 399.680000 154.460000 400.520000 ;
      RECT 151.900000 399.680000 153.080000 400.520000 ;
      RECT 150.520000 399.680000 151.240000 400.520000 ;
      RECT 149.140000 399.680000 149.860000 400.520000 ;
      RECT 147.300000 399.680000 148.480000 400.520000 ;
      RECT 145.920000 399.680000 146.640000 400.520000 ;
      RECT 144.540000 399.680000 145.260000 400.520000 ;
      RECT 143.160000 399.680000 143.880000 400.520000 ;
      RECT 141.320000 399.680000 142.500000 400.520000 ;
      RECT 139.940000 399.680000 140.660000 400.520000 ;
      RECT 138.560000 399.680000 139.280000 400.520000 ;
      RECT 136.720000 399.680000 137.900000 400.520000 ;
      RECT 135.340000 399.680000 136.060000 400.520000 ;
      RECT 133.960000 399.680000 134.680000 400.520000 ;
      RECT 132.120000 399.680000 133.300000 400.520000 ;
      RECT 130.740000 399.680000 131.460000 400.520000 ;
      RECT 129.360000 399.680000 130.080000 400.520000 ;
      RECT 127.520000 399.680000 128.700000 400.520000 ;
      RECT 126.140000 399.680000 126.860000 400.520000 ;
      RECT 124.760000 399.680000 125.480000 400.520000 ;
      RECT 122.920000 399.680000 124.100000 400.520000 ;
      RECT 121.540000 399.680000 122.260000 400.520000 ;
      RECT 120.160000 399.680000 120.880000 400.520000 ;
      RECT 118.320000 399.680000 119.500000 400.520000 ;
      RECT 116.940000 399.680000 117.660000 400.520000 ;
      RECT 115.560000 399.680000 116.280000 400.520000 ;
      RECT 113.720000 399.680000 114.900000 400.520000 ;
      RECT 112.340000 399.680000 113.060000 400.520000 ;
      RECT 110.960000 399.680000 111.680000 400.520000 ;
      RECT 109.120000 399.680000 110.300000 400.520000 ;
      RECT 107.740000 399.680000 108.460000 400.520000 ;
      RECT 106.360000 399.680000 107.080000 400.520000 ;
      RECT 104.520000 399.680000 105.700000 400.520000 ;
      RECT 103.140000 399.680000 103.860000 400.520000 ;
      RECT 101.760000 399.680000 102.480000 400.520000 ;
      RECT 99.920000 399.680000 101.100000 400.520000 ;
      RECT 98.540000 399.680000 99.260000 400.520000 ;
      RECT 97.160000 399.680000 97.880000 400.520000 ;
      RECT 95.780000 399.680000 96.500000 400.520000 ;
      RECT 93.940000 399.680000 95.120000 400.520000 ;
      RECT 92.560000 399.680000 93.280000 400.520000 ;
      RECT 91.180000 399.680000 91.900000 400.520000 ;
      RECT 89.340000 399.680000 90.520000 400.520000 ;
      RECT 87.960000 399.680000 88.680000 400.520000 ;
      RECT 86.580000 399.680000 87.300000 400.520000 ;
      RECT 84.740000 399.680000 85.920000 400.520000 ;
      RECT 83.360000 399.680000 84.080000 400.520000 ;
      RECT 81.980000 399.680000 82.700000 400.520000 ;
      RECT 80.140000 399.680000 81.320000 400.520000 ;
      RECT 78.760000 399.680000 79.480000 400.520000 ;
      RECT 77.380000 399.680000 78.100000 400.520000 ;
      RECT 75.540000 399.680000 76.720000 400.520000 ;
      RECT 74.160000 399.680000 74.880000 400.520000 ;
      RECT 72.780000 399.680000 73.500000 400.520000 ;
      RECT 70.940000 399.680000 72.120000 400.520000 ;
      RECT 69.560000 399.680000 70.280000 400.520000 ;
      RECT 68.180000 399.680000 68.900000 400.520000 ;
      RECT 66.340000 399.680000 67.520000 400.520000 ;
      RECT 64.960000 399.680000 65.680000 400.520000 ;
      RECT 63.580000 399.680000 64.300000 400.520000 ;
      RECT 61.740000 399.680000 62.920000 400.520000 ;
      RECT 60.360000 399.680000 61.080000 400.520000 ;
      RECT 58.980000 399.680000 59.700000 400.520000 ;
      RECT 57.140000 399.680000 58.320000 400.520000 ;
      RECT 55.760000 399.680000 56.480000 400.520000 ;
      RECT 54.380000 399.680000 55.100000 400.520000 ;
      RECT 53.000000 399.680000 53.720000 400.520000 ;
      RECT 51.160000 399.680000 52.340000 400.520000 ;
      RECT 49.780000 399.680000 50.500000 400.520000 ;
      RECT 48.400000 399.680000 49.120000 400.520000 ;
      RECT 46.560000 399.680000 47.740000 400.520000 ;
      RECT 45.180000 399.680000 45.900000 400.520000 ;
      RECT 43.800000 399.680000 44.520000 400.520000 ;
      RECT 41.960000 399.680000 43.140000 400.520000 ;
      RECT 40.580000 399.680000 41.300000 400.520000 ;
      RECT 39.200000 399.680000 39.920000 400.520000 ;
      RECT 37.360000 399.680000 38.540000 400.520000 ;
      RECT 35.980000 399.680000 36.700000 400.520000 ;
      RECT 34.600000 399.680000 35.320000 400.520000 ;
      RECT 32.760000 399.680000 33.940000 400.520000 ;
      RECT 31.380000 399.680000 32.100000 400.520000 ;
      RECT 30.000000 399.680000 30.720000 400.520000 ;
      RECT 28.160000 399.680000 29.340000 400.520000 ;
      RECT 26.780000 399.680000 27.500000 400.520000 ;
      RECT 25.400000 399.680000 26.120000 400.520000 ;
      RECT 23.560000 399.680000 24.740000 400.520000 ;
      RECT 22.180000 399.680000 22.900000 400.520000 ;
      RECT 20.800000 399.680000 21.520000 400.520000 ;
      RECT 18.960000 399.680000 20.140000 400.520000 ;
      RECT 17.580000 399.680000 18.300000 400.520000 ;
      RECT 16.200000 399.680000 16.920000 400.520000 ;
      RECT 14.360000 399.680000 15.540000 400.520000 ;
      RECT 12.980000 399.680000 13.700000 400.520000 ;
      RECT 11.600000 399.680000 12.320000 400.520000 ;
      RECT 9.760000 399.680000 10.940000 400.520000 ;
      RECT 8.380000 399.680000 9.100000 400.520000 ;
      RECT 7.000000 399.680000 7.720000 400.520000 ;
      RECT 5.620000 399.680000 6.340000 400.520000 ;
      RECT 0.000000 399.680000 4.960000 400.520000 ;
      RECT 0.000000 0.840000 200.100000 399.680000 ;
      RECT 194.680000 0.000000 200.100000 0.840000 ;
      RECT 193.300000 0.000000 194.020000 0.840000 ;
      RECT 191.920000 0.000000 192.640000 0.840000 ;
      RECT 190.540000 0.000000 191.260000 0.840000 ;
      RECT 188.700000 0.000000 189.880000 0.840000 ;
      RECT 187.320000 0.000000 188.040000 0.840000 ;
      RECT 185.940000 0.000000 186.660000 0.840000 ;
      RECT 184.100000 0.000000 185.280000 0.840000 ;
      RECT 182.720000 0.000000 183.440000 0.840000 ;
      RECT 181.340000 0.000000 182.060000 0.840000 ;
      RECT 179.500000 0.000000 180.680000 0.840000 ;
      RECT 178.120000 0.000000 178.840000 0.840000 ;
      RECT 176.740000 0.000000 177.460000 0.840000 ;
      RECT 174.900000 0.000000 176.080000 0.840000 ;
      RECT 173.520000 0.000000 174.240000 0.840000 ;
      RECT 172.140000 0.000000 172.860000 0.840000 ;
      RECT 170.300000 0.000000 171.480000 0.840000 ;
      RECT 168.920000 0.000000 169.640000 0.840000 ;
      RECT 167.540000 0.000000 168.260000 0.840000 ;
      RECT 165.700000 0.000000 166.880000 0.840000 ;
      RECT 164.320000 0.000000 165.040000 0.840000 ;
      RECT 162.940000 0.000000 163.660000 0.840000 ;
      RECT 161.100000 0.000000 162.280000 0.840000 ;
      RECT 159.720000 0.000000 160.440000 0.840000 ;
      RECT 158.340000 0.000000 159.060000 0.840000 ;
      RECT 156.500000 0.000000 157.680000 0.840000 ;
      RECT 155.120000 0.000000 155.840000 0.840000 ;
      RECT 153.740000 0.000000 154.460000 0.840000 ;
      RECT 151.900000 0.000000 153.080000 0.840000 ;
      RECT 150.520000 0.000000 151.240000 0.840000 ;
      RECT 149.140000 0.000000 149.860000 0.840000 ;
      RECT 147.300000 0.000000 148.480000 0.840000 ;
      RECT 145.920000 0.000000 146.640000 0.840000 ;
      RECT 144.540000 0.000000 145.260000 0.840000 ;
      RECT 143.160000 0.000000 143.880000 0.840000 ;
      RECT 141.320000 0.000000 142.500000 0.840000 ;
      RECT 139.940000 0.000000 140.660000 0.840000 ;
      RECT 138.560000 0.000000 139.280000 0.840000 ;
      RECT 136.720000 0.000000 137.900000 0.840000 ;
      RECT 135.340000 0.000000 136.060000 0.840000 ;
      RECT 133.960000 0.000000 134.680000 0.840000 ;
      RECT 132.120000 0.000000 133.300000 0.840000 ;
      RECT 130.740000 0.000000 131.460000 0.840000 ;
      RECT 129.360000 0.000000 130.080000 0.840000 ;
      RECT 127.520000 0.000000 128.700000 0.840000 ;
      RECT 126.140000 0.000000 126.860000 0.840000 ;
      RECT 124.760000 0.000000 125.480000 0.840000 ;
      RECT 122.920000 0.000000 124.100000 0.840000 ;
      RECT 121.540000 0.000000 122.260000 0.840000 ;
      RECT 120.160000 0.000000 120.880000 0.840000 ;
      RECT 118.320000 0.000000 119.500000 0.840000 ;
      RECT 116.940000 0.000000 117.660000 0.840000 ;
      RECT 115.560000 0.000000 116.280000 0.840000 ;
      RECT 113.720000 0.000000 114.900000 0.840000 ;
      RECT 112.340000 0.000000 113.060000 0.840000 ;
      RECT 110.960000 0.000000 111.680000 0.840000 ;
      RECT 109.120000 0.000000 110.300000 0.840000 ;
      RECT 107.740000 0.000000 108.460000 0.840000 ;
      RECT 106.360000 0.000000 107.080000 0.840000 ;
      RECT 104.520000 0.000000 105.700000 0.840000 ;
      RECT 103.140000 0.000000 103.860000 0.840000 ;
      RECT 101.760000 0.000000 102.480000 0.840000 ;
      RECT 99.920000 0.000000 101.100000 0.840000 ;
      RECT 98.540000 0.000000 99.260000 0.840000 ;
      RECT 97.160000 0.000000 97.880000 0.840000 ;
      RECT 95.780000 0.000000 96.500000 0.840000 ;
      RECT 93.940000 0.000000 95.120000 0.840000 ;
      RECT 92.560000 0.000000 93.280000 0.840000 ;
      RECT 91.180000 0.000000 91.900000 0.840000 ;
      RECT 89.340000 0.000000 90.520000 0.840000 ;
      RECT 87.960000 0.000000 88.680000 0.840000 ;
      RECT 86.580000 0.000000 87.300000 0.840000 ;
      RECT 84.740000 0.000000 85.920000 0.840000 ;
      RECT 83.360000 0.000000 84.080000 0.840000 ;
      RECT 81.980000 0.000000 82.700000 0.840000 ;
      RECT 80.140000 0.000000 81.320000 0.840000 ;
      RECT 78.760000 0.000000 79.480000 0.840000 ;
      RECT 77.380000 0.000000 78.100000 0.840000 ;
      RECT 75.540000 0.000000 76.720000 0.840000 ;
      RECT 74.160000 0.000000 74.880000 0.840000 ;
      RECT 72.780000 0.000000 73.500000 0.840000 ;
      RECT 70.940000 0.000000 72.120000 0.840000 ;
      RECT 69.560000 0.000000 70.280000 0.840000 ;
      RECT 68.180000 0.000000 68.900000 0.840000 ;
      RECT 66.340000 0.000000 67.520000 0.840000 ;
      RECT 64.960000 0.000000 65.680000 0.840000 ;
      RECT 63.580000 0.000000 64.300000 0.840000 ;
      RECT 61.740000 0.000000 62.920000 0.840000 ;
      RECT 60.360000 0.000000 61.080000 0.840000 ;
      RECT 58.980000 0.000000 59.700000 0.840000 ;
      RECT 57.140000 0.000000 58.320000 0.840000 ;
      RECT 55.760000 0.000000 56.480000 0.840000 ;
      RECT 54.380000 0.000000 55.100000 0.840000 ;
      RECT 53.000000 0.000000 53.720000 0.840000 ;
      RECT 51.160000 0.000000 52.340000 0.840000 ;
      RECT 49.780000 0.000000 50.500000 0.840000 ;
      RECT 48.400000 0.000000 49.120000 0.840000 ;
      RECT 46.560000 0.000000 47.740000 0.840000 ;
      RECT 45.180000 0.000000 45.900000 0.840000 ;
      RECT 43.800000 0.000000 44.520000 0.840000 ;
      RECT 41.960000 0.000000 43.140000 0.840000 ;
      RECT 40.580000 0.000000 41.300000 0.840000 ;
      RECT 39.200000 0.000000 39.920000 0.840000 ;
      RECT 37.360000 0.000000 38.540000 0.840000 ;
      RECT 35.980000 0.000000 36.700000 0.840000 ;
      RECT 34.600000 0.000000 35.320000 0.840000 ;
      RECT 32.760000 0.000000 33.940000 0.840000 ;
      RECT 31.380000 0.000000 32.100000 0.840000 ;
      RECT 30.000000 0.000000 30.720000 0.840000 ;
      RECT 28.160000 0.000000 29.340000 0.840000 ;
      RECT 26.780000 0.000000 27.500000 0.840000 ;
      RECT 25.400000 0.000000 26.120000 0.840000 ;
      RECT 23.560000 0.000000 24.740000 0.840000 ;
      RECT 22.180000 0.000000 22.900000 0.840000 ;
      RECT 20.800000 0.000000 21.520000 0.840000 ;
      RECT 18.960000 0.000000 20.140000 0.840000 ;
      RECT 17.580000 0.000000 18.300000 0.840000 ;
      RECT 16.200000 0.000000 16.920000 0.840000 ;
      RECT 14.360000 0.000000 15.540000 0.840000 ;
      RECT 12.980000 0.000000 13.700000 0.840000 ;
      RECT 11.600000 0.000000 12.320000 0.840000 ;
      RECT 9.760000 0.000000 10.940000 0.840000 ;
      RECT 8.380000 0.000000 9.100000 0.840000 ;
      RECT 7.000000 0.000000 7.720000 0.840000 ;
      RECT 5.620000 0.000000 6.340000 0.840000 ;
      RECT 0.000000 0.000000 4.960000 0.840000 ;
    LAYER met3 ;
      RECT 0.000000 399.090000 200.100000 400.520000 ;
      RECT 0.000000 394.940000 200.100000 395.490000 ;
      RECT 1.000000 394.600000 199.100000 394.940000 ;
      RECT 199.370000 393.520000 200.100000 393.960000 ;
      RECT 186.560000 393.520000 197.570000 394.600000 ;
      RECT 141.560000 393.520000 184.760000 394.600000 ;
      RECT 96.560000 393.520000 139.760000 394.600000 ;
      RECT 51.560000 393.520000 94.760000 394.600000 ;
      RECT 6.560000 393.520000 49.760000 394.600000 ;
      RECT 2.530000 393.520000 4.595000 394.600000 ;
      RECT 0.000000 393.520000 0.730000 393.960000 ;
      RECT 0.000000 393.110000 200.100000 393.520000 ;
      RECT 1.000000 392.130000 199.100000 393.110000 ;
      RECT 0.000000 391.890000 200.100000 392.130000 ;
      RECT 1.000000 391.880000 199.100000 391.890000 ;
      RECT 197.570000 390.910000 199.100000 391.880000 ;
      RECT 1.000000 390.910000 2.530000 391.880000 ;
      RECT 197.570000 390.800000 200.100000 390.910000 ;
      RECT 188.560000 390.800000 195.770000 391.880000 ;
      RECT 143.560000 390.800000 186.760000 391.880000 ;
      RECT 98.560000 390.800000 141.760000 391.880000 ;
      RECT 53.560000 390.800000 96.760000 391.880000 ;
      RECT 8.560000 390.800000 51.760000 391.880000 ;
      RECT 4.330000 390.800000 6.760000 391.880000 ;
      RECT 0.000000 390.800000 2.530000 390.910000 ;
      RECT 0.000000 390.060000 200.100000 390.800000 ;
      RECT 1.000000 389.160000 199.100000 390.060000 ;
      RECT 199.370000 388.840000 200.100000 389.080000 ;
      RECT 0.000000 388.840000 0.730000 389.080000 ;
      RECT 186.560000 388.080000 197.570000 389.160000 ;
      RECT 141.560000 388.080000 184.760000 389.160000 ;
      RECT 96.560000 388.080000 139.760000 389.160000 ;
      RECT 51.560000 388.080000 94.760000 389.160000 ;
      RECT 6.560000 388.080000 49.760000 389.160000 ;
      RECT 2.530000 388.080000 4.595000 389.160000 ;
      RECT 1.000000 387.860000 199.100000 388.080000 ;
      RECT 0.000000 387.010000 200.100000 387.860000 ;
      RECT 1.000000 386.440000 199.100000 387.010000 ;
      RECT 197.570000 386.030000 199.100000 386.440000 ;
      RECT 1.000000 386.030000 2.530000 386.440000 ;
      RECT 197.570000 385.790000 200.100000 386.030000 ;
      RECT 0.000000 385.790000 2.530000 386.030000 ;
      RECT 197.570000 385.360000 199.100000 385.790000 ;
      RECT 188.560000 385.360000 195.770000 386.440000 ;
      RECT 143.560000 385.360000 186.760000 386.440000 ;
      RECT 98.560000 385.360000 141.760000 386.440000 ;
      RECT 53.560000 385.360000 96.760000 386.440000 ;
      RECT 8.560000 385.360000 51.760000 386.440000 ;
      RECT 4.330000 385.360000 6.760000 386.440000 ;
      RECT 1.000000 385.360000 2.530000 385.790000 ;
      RECT 1.000000 384.810000 199.100000 385.360000 ;
      RECT 0.000000 383.960000 200.100000 384.810000 ;
      RECT 1.000000 383.720000 199.100000 383.960000 ;
      RECT 199.370000 382.740000 200.100000 382.980000 ;
      RECT 0.000000 382.740000 0.730000 382.980000 ;
      RECT 186.560000 382.640000 197.570000 383.720000 ;
      RECT 141.560000 382.640000 184.760000 383.720000 ;
      RECT 96.560000 382.640000 139.760000 383.720000 ;
      RECT 51.560000 382.640000 94.760000 383.720000 ;
      RECT 6.560000 382.640000 49.760000 383.720000 ;
      RECT 2.530000 382.640000 4.595000 383.720000 ;
      RECT 1.000000 381.760000 199.100000 382.640000 ;
      RECT 0.000000 381.520000 200.100000 381.760000 ;
      RECT 1.000000 381.000000 199.100000 381.520000 ;
      RECT 197.570000 380.540000 199.100000 381.000000 ;
      RECT 1.000000 380.540000 2.530000 381.000000 ;
      RECT 197.570000 379.920000 200.100000 380.540000 ;
      RECT 188.560000 379.920000 195.770000 381.000000 ;
      RECT 143.560000 379.920000 186.760000 381.000000 ;
      RECT 98.560000 379.920000 141.760000 381.000000 ;
      RECT 53.560000 379.920000 96.760000 381.000000 ;
      RECT 8.560000 379.920000 51.760000 381.000000 ;
      RECT 4.330000 379.920000 6.760000 381.000000 ;
      RECT 0.000000 379.920000 2.530000 380.540000 ;
      RECT 0.000000 379.690000 200.100000 379.920000 ;
      RECT 1.000000 378.710000 199.100000 379.690000 ;
      RECT 0.000000 378.470000 200.100000 378.710000 ;
      RECT 1.000000 378.280000 199.100000 378.470000 ;
      RECT 199.370000 377.200000 200.100000 377.490000 ;
      RECT 186.560000 377.200000 197.570000 378.280000 ;
      RECT 141.560000 377.200000 184.760000 378.280000 ;
      RECT 96.560000 377.200000 139.760000 378.280000 ;
      RECT 51.560000 377.200000 94.760000 378.280000 ;
      RECT 6.560000 377.200000 49.760000 378.280000 ;
      RECT 2.530000 377.200000 4.595000 378.280000 ;
      RECT 0.000000 377.200000 0.730000 377.490000 ;
      RECT 0.000000 376.640000 200.100000 377.200000 ;
      RECT 1.000000 375.660000 199.100000 376.640000 ;
      RECT 0.000000 375.560000 200.100000 375.660000 ;
      RECT 197.570000 375.420000 200.100000 375.560000 ;
      RECT 0.000000 375.420000 2.530000 375.560000 ;
      RECT 197.570000 374.480000 199.100000 375.420000 ;
      RECT 188.560000 374.480000 195.770000 375.560000 ;
      RECT 143.560000 374.480000 186.760000 375.560000 ;
      RECT 98.560000 374.480000 141.760000 375.560000 ;
      RECT 53.560000 374.480000 96.760000 375.560000 ;
      RECT 8.560000 374.480000 51.760000 375.560000 ;
      RECT 4.330000 374.480000 6.760000 375.560000 ;
      RECT 1.000000 374.480000 2.530000 375.420000 ;
      RECT 1.000000 374.440000 199.100000 374.480000 ;
      RECT 0.000000 373.590000 200.100000 374.440000 ;
      RECT 1.000000 372.840000 199.100000 373.590000 ;
      RECT 199.370000 372.370000 200.100000 372.610000 ;
      RECT 0.000000 372.370000 0.730000 372.610000 ;
      RECT 186.560000 371.760000 197.570000 372.840000 ;
      RECT 141.560000 371.760000 184.760000 372.840000 ;
      RECT 96.560000 371.760000 139.760000 372.840000 ;
      RECT 51.560000 371.760000 94.760000 372.840000 ;
      RECT 6.560000 371.760000 49.760000 372.840000 ;
      RECT 2.530000 371.760000 4.595000 372.840000 ;
      RECT 1.000000 371.390000 199.100000 371.760000 ;
      RECT 0.000000 370.540000 200.100000 371.390000 ;
      RECT 1.000000 370.120000 199.100000 370.540000 ;
      RECT 197.570000 369.560000 199.100000 370.120000 ;
      RECT 1.000000 369.560000 2.530000 370.120000 ;
      RECT 197.570000 369.320000 200.100000 369.560000 ;
      RECT 0.000000 369.320000 2.530000 369.560000 ;
      RECT 197.570000 369.040000 199.100000 369.320000 ;
      RECT 188.560000 369.040000 195.770000 370.120000 ;
      RECT 143.560000 369.040000 186.760000 370.120000 ;
      RECT 98.560000 369.040000 141.760000 370.120000 ;
      RECT 53.560000 369.040000 96.760000 370.120000 ;
      RECT 8.560000 369.040000 51.760000 370.120000 ;
      RECT 4.330000 369.040000 6.760000 370.120000 ;
      RECT 1.000000 369.040000 2.530000 369.320000 ;
      RECT 1.000000 368.340000 199.100000 369.040000 ;
      RECT 0.000000 368.100000 200.100000 368.340000 ;
      RECT 1.000000 367.400000 199.100000 368.100000 ;
      RECT 199.370000 366.320000 200.100000 367.120000 ;
      RECT 186.560000 366.320000 197.570000 367.400000 ;
      RECT 141.560000 366.320000 184.760000 367.400000 ;
      RECT 96.560000 366.320000 139.760000 367.400000 ;
      RECT 51.560000 366.320000 94.760000 367.400000 ;
      RECT 6.560000 366.320000 49.760000 367.400000 ;
      RECT 2.530000 366.320000 4.595000 367.400000 ;
      RECT 0.000000 366.320000 0.730000 367.120000 ;
      RECT 0.000000 366.270000 200.100000 366.320000 ;
      RECT 1.000000 365.290000 199.100000 366.270000 ;
      RECT 0.000000 365.050000 200.100000 365.290000 ;
      RECT 1.000000 364.680000 199.100000 365.050000 ;
      RECT 197.570000 364.070000 199.100000 364.680000 ;
      RECT 1.000000 364.070000 2.530000 364.680000 ;
      RECT 197.570000 363.600000 200.100000 364.070000 ;
      RECT 188.560000 363.600000 195.770000 364.680000 ;
      RECT 143.560000 363.600000 186.760000 364.680000 ;
      RECT 98.560000 363.600000 141.760000 364.680000 ;
      RECT 53.560000 363.600000 96.760000 364.680000 ;
      RECT 8.560000 363.600000 51.760000 364.680000 ;
      RECT 4.330000 363.600000 6.760000 364.680000 ;
      RECT 0.000000 363.600000 2.530000 364.070000 ;
      RECT 0.000000 363.220000 200.100000 363.600000 ;
      RECT 1.000000 362.240000 199.100000 363.220000 ;
      RECT 0.000000 362.000000 200.100000 362.240000 ;
      RECT 1.000000 361.960000 199.100000 362.000000 ;
      RECT 199.370000 360.880000 200.100000 361.020000 ;
      RECT 186.560000 360.880000 197.570000 361.960000 ;
      RECT 141.560000 360.880000 184.760000 361.960000 ;
      RECT 96.560000 360.880000 139.760000 361.960000 ;
      RECT 51.560000 360.880000 94.760000 361.960000 ;
      RECT 6.560000 360.880000 49.760000 361.960000 ;
      RECT 2.530000 360.880000 4.595000 361.960000 ;
      RECT 0.000000 360.880000 0.730000 361.020000 ;
      RECT 0.000000 360.170000 200.100000 360.880000 ;
      RECT 1.000000 359.240000 199.100000 360.170000 ;
      RECT 197.570000 359.190000 199.100000 359.240000 ;
      RECT 1.000000 359.190000 2.530000 359.240000 ;
      RECT 197.570000 358.950000 200.100000 359.190000 ;
      RECT 0.000000 358.950000 2.530000 359.190000 ;
      RECT 197.570000 358.160000 199.100000 358.950000 ;
      RECT 188.560000 358.160000 195.770000 359.240000 ;
      RECT 143.560000 358.160000 186.760000 359.240000 ;
      RECT 98.560000 358.160000 141.760000 359.240000 ;
      RECT 53.560000 358.160000 96.760000 359.240000 ;
      RECT 8.560000 358.160000 51.760000 359.240000 ;
      RECT 4.330000 358.160000 6.760000 359.240000 ;
      RECT 1.000000 358.160000 2.530000 358.950000 ;
      RECT 1.000000 357.970000 199.100000 358.160000 ;
      RECT 0.000000 357.120000 200.100000 357.970000 ;
      RECT 1.000000 356.520000 199.100000 357.120000 ;
      RECT 199.370000 355.900000 200.100000 356.140000 ;
      RECT 0.000000 355.900000 0.730000 356.140000 ;
      RECT 186.560000 355.440000 197.570000 356.520000 ;
      RECT 141.560000 355.440000 184.760000 356.520000 ;
      RECT 96.560000 355.440000 139.760000 356.520000 ;
      RECT 51.560000 355.440000 94.760000 356.520000 ;
      RECT 6.560000 355.440000 49.760000 356.520000 ;
      RECT 2.530000 355.440000 4.595000 356.520000 ;
      RECT 1.000000 354.920000 199.100000 355.440000 ;
      RECT 0.000000 354.680000 200.100000 354.920000 ;
      RECT 1.000000 353.800000 199.100000 354.680000 ;
      RECT 197.570000 353.700000 199.100000 353.800000 ;
      RECT 1.000000 353.700000 2.530000 353.800000 ;
      RECT 197.570000 352.850000 200.100000 353.700000 ;
      RECT 0.000000 352.850000 2.530000 353.700000 ;
      RECT 197.570000 352.720000 199.100000 352.850000 ;
      RECT 188.560000 352.720000 195.770000 353.800000 ;
      RECT 143.560000 352.720000 186.760000 353.800000 ;
      RECT 98.560000 352.720000 141.760000 353.800000 ;
      RECT 53.560000 352.720000 96.760000 353.800000 ;
      RECT 8.560000 352.720000 51.760000 353.800000 ;
      RECT 4.330000 352.720000 6.760000 353.800000 ;
      RECT 1.000000 352.720000 2.530000 352.850000 ;
      RECT 1.000000 351.870000 199.100000 352.720000 ;
      RECT 0.000000 351.630000 200.100000 351.870000 ;
      RECT 1.000000 351.080000 199.100000 351.630000 ;
      RECT 199.370000 350.000000 200.100000 350.650000 ;
      RECT 186.560000 350.000000 197.570000 351.080000 ;
      RECT 141.560000 350.000000 184.760000 351.080000 ;
      RECT 96.560000 350.000000 139.760000 351.080000 ;
      RECT 51.560000 350.000000 94.760000 351.080000 ;
      RECT 6.560000 350.000000 49.760000 351.080000 ;
      RECT 2.530000 350.000000 4.595000 351.080000 ;
      RECT 0.000000 350.000000 0.730000 350.650000 ;
      RECT 0.000000 349.800000 200.100000 350.000000 ;
      RECT 1.000000 348.820000 199.100000 349.800000 ;
      RECT 0.000000 348.580000 200.100000 348.820000 ;
      RECT 1.000000 348.360000 199.100000 348.580000 ;
      RECT 197.570000 347.600000 199.100000 348.360000 ;
      RECT 1.000000 347.600000 2.530000 348.360000 ;
      RECT 197.570000 347.280000 200.100000 347.600000 ;
      RECT 188.560000 347.280000 195.770000 348.360000 ;
      RECT 143.560000 347.280000 186.760000 348.360000 ;
      RECT 98.560000 347.280000 141.760000 348.360000 ;
      RECT 53.560000 347.280000 96.760000 348.360000 ;
      RECT 8.560000 347.280000 51.760000 348.360000 ;
      RECT 4.330000 347.280000 6.760000 348.360000 ;
      RECT 0.000000 347.280000 2.530000 347.600000 ;
      RECT 0.000000 346.750000 200.100000 347.280000 ;
      RECT 1.000000 345.770000 199.100000 346.750000 ;
      RECT 0.000000 345.640000 200.100000 345.770000 ;
      RECT 199.370000 345.530000 200.100000 345.640000 ;
      RECT 0.000000 345.530000 0.730000 345.640000 ;
      RECT 186.560000 344.560000 197.570000 345.640000 ;
      RECT 141.560000 344.560000 184.760000 345.640000 ;
      RECT 96.560000 344.560000 139.760000 345.640000 ;
      RECT 51.560000 344.560000 94.760000 345.640000 ;
      RECT 6.560000 344.560000 49.760000 345.640000 ;
      RECT 2.530000 344.560000 4.595000 345.640000 ;
      RECT 1.000000 344.550000 199.100000 344.560000 ;
      RECT 0.000000 344.310000 200.100000 344.550000 ;
      RECT 1.000000 343.330000 199.100000 344.310000 ;
      RECT 0.000000 342.920000 200.100000 343.330000 ;
      RECT 197.570000 342.480000 200.100000 342.920000 ;
      RECT 0.000000 342.480000 2.530000 342.920000 ;
      RECT 197.570000 341.840000 199.100000 342.480000 ;
      RECT 188.560000 341.840000 195.770000 342.920000 ;
      RECT 143.560000 341.840000 186.760000 342.920000 ;
      RECT 98.560000 341.840000 141.760000 342.920000 ;
      RECT 53.560000 341.840000 96.760000 342.920000 ;
      RECT 8.560000 341.840000 51.760000 342.920000 ;
      RECT 4.330000 341.840000 6.760000 342.920000 ;
      RECT 1.000000 341.840000 2.530000 342.480000 ;
      RECT 1.000000 341.500000 199.100000 341.840000 ;
      RECT 0.000000 341.260000 200.100000 341.500000 ;
      RECT 1.000000 340.280000 199.100000 341.260000 ;
      RECT 0.000000 340.200000 200.100000 340.280000 ;
      RECT 199.370000 339.430000 200.100000 340.200000 ;
      RECT 0.000000 339.430000 0.730000 340.200000 ;
      RECT 186.560000 339.120000 197.570000 340.200000 ;
      RECT 141.560000 339.120000 184.760000 340.200000 ;
      RECT 96.560000 339.120000 139.760000 340.200000 ;
      RECT 51.560000 339.120000 94.760000 340.200000 ;
      RECT 6.560000 339.120000 49.760000 340.200000 ;
      RECT 2.530000 339.120000 4.595000 340.200000 ;
      RECT 1.000000 338.450000 199.100000 339.120000 ;
      RECT 0.000000 338.210000 200.100000 338.450000 ;
      RECT 1.000000 337.480000 199.100000 338.210000 ;
      RECT 197.570000 337.230000 199.100000 337.480000 ;
      RECT 1.000000 337.230000 2.530000 337.480000 ;
      RECT 197.570000 336.400000 200.100000 337.230000 ;
      RECT 188.560000 336.400000 195.770000 337.480000 ;
      RECT 143.560000 336.400000 186.760000 337.480000 ;
      RECT 98.560000 336.400000 141.760000 337.480000 ;
      RECT 53.560000 336.400000 96.760000 337.480000 ;
      RECT 8.560000 336.400000 51.760000 337.480000 ;
      RECT 4.330000 336.400000 6.760000 337.480000 ;
      RECT 0.000000 336.400000 2.530000 337.230000 ;
      RECT 0.000000 336.380000 200.100000 336.400000 ;
      RECT 1.000000 335.400000 199.100000 336.380000 ;
      RECT 0.000000 335.160000 200.100000 335.400000 ;
      RECT 1.000000 334.760000 199.100000 335.160000 ;
      RECT 199.370000 333.680000 200.100000 334.180000 ;
      RECT 186.560000 333.680000 197.570000 334.760000 ;
      RECT 141.560000 333.680000 184.760000 334.760000 ;
      RECT 96.560000 333.680000 139.760000 334.760000 ;
      RECT 51.560000 333.680000 94.760000 334.760000 ;
      RECT 6.560000 333.680000 49.760000 334.760000 ;
      RECT 2.530000 333.680000 4.595000 334.760000 ;
      RECT 0.000000 333.680000 0.730000 334.180000 ;
      RECT 0.000000 333.330000 200.100000 333.680000 ;
      RECT 1.000000 332.350000 199.100000 333.330000 ;
      RECT 0.000000 332.110000 200.100000 332.350000 ;
      RECT 1.000000 332.040000 199.100000 332.110000 ;
      RECT 197.570000 331.130000 199.100000 332.040000 ;
      RECT 1.000000 331.130000 2.530000 332.040000 ;
      RECT 197.570000 330.960000 200.100000 331.130000 ;
      RECT 188.560000 330.960000 195.770000 332.040000 ;
      RECT 143.560000 330.960000 186.760000 332.040000 ;
      RECT 98.560000 330.960000 141.760000 332.040000 ;
      RECT 53.560000 330.960000 96.760000 332.040000 ;
      RECT 8.560000 330.960000 51.760000 332.040000 ;
      RECT 4.330000 330.960000 6.760000 332.040000 ;
      RECT 0.000000 330.960000 2.530000 331.130000 ;
      RECT 0.000000 330.890000 200.100000 330.960000 ;
      RECT 1.000000 329.910000 199.100000 330.890000 ;
      RECT 0.000000 329.320000 200.100000 329.910000 ;
      RECT 199.370000 329.060000 200.100000 329.320000 ;
      RECT 0.000000 329.060000 0.730000 329.320000 ;
      RECT 186.560000 328.240000 197.570000 329.320000 ;
      RECT 141.560000 328.240000 184.760000 329.320000 ;
      RECT 96.560000 328.240000 139.760000 329.320000 ;
      RECT 51.560000 328.240000 94.760000 329.320000 ;
      RECT 6.560000 328.240000 49.760000 329.320000 ;
      RECT 2.530000 328.240000 4.595000 329.320000 ;
      RECT 1.000000 328.080000 199.100000 328.240000 ;
      RECT 0.000000 327.840000 200.100000 328.080000 ;
      RECT 1.000000 326.860000 199.100000 327.840000 ;
      RECT 0.000000 326.600000 200.100000 326.860000 ;
      RECT 197.570000 326.010000 200.100000 326.600000 ;
      RECT 0.000000 326.010000 2.530000 326.600000 ;
      RECT 197.570000 325.520000 199.100000 326.010000 ;
      RECT 188.560000 325.520000 195.770000 326.600000 ;
      RECT 143.560000 325.520000 186.760000 326.600000 ;
      RECT 98.560000 325.520000 141.760000 326.600000 ;
      RECT 53.560000 325.520000 96.760000 326.600000 ;
      RECT 8.560000 325.520000 51.760000 326.600000 ;
      RECT 4.330000 325.520000 6.760000 326.600000 ;
      RECT 1.000000 325.520000 2.530000 326.010000 ;
      RECT 1.000000 325.030000 199.100000 325.520000 ;
      RECT 0.000000 324.790000 200.100000 325.030000 ;
      RECT 1.000000 323.880000 199.100000 324.790000 ;
      RECT 199.370000 322.960000 200.100000 323.810000 ;
      RECT 0.000000 322.960000 0.730000 323.810000 ;
      RECT 186.560000 322.800000 197.570000 323.880000 ;
      RECT 141.560000 322.800000 184.760000 323.880000 ;
      RECT 96.560000 322.800000 139.760000 323.880000 ;
      RECT 51.560000 322.800000 94.760000 323.880000 ;
      RECT 6.560000 322.800000 49.760000 323.880000 ;
      RECT 2.530000 322.800000 4.595000 323.880000 ;
      RECT 1.000000 321.980000 199.100000 322.800000 ;
      RECT 0.000000 321.740000 200.100000 321.980000 ;
      RECT 1.000000 321.160000 199.100000 321.740000 ;
      RECT 197.570000 320.760000 199.100000 321.160000 ;
      RECT 1.000000 320.760000 2.530000 321.160000 ;
      RECT 197.570000 320.080000 200.100000 320.760000 ;
      RECT 188.560000 320.080000 195.770000 321.160000 ;
      RECT 143.560000 320.080000 186.760000 321.160000 ;
      RECT 98.560000 320.080000 141.760000 321.160000 ;
      RECT 53.560000 320.080000 96.760000 321.160000 ;
      RECT 8.560000 320.080000 51.760000 321.160000 ;
      RECT 4.330000 320.080000 6.760000 321.160000 ;
      RECT 0.000000 320.080000 2.530000 320.760000 ;
      RECT 0.000000 319.910000 200.100000 320.080000 ;
      RECT 1.000000 318.930000 199.100000 319.910000 ;
      RECT 0.000000 318.690000 200.100000 318.930000 ;
      RECT 1.000000 318.440000 199.100000 318.690000 ;
      RECT 199.370000 317.470000 200.100000 317.710000 ;
      RECT 0.000000 317.470000 0.730000 317.710000 ;
      RECT 186.560000 317.360000 197.570000 318.440000 ;
      RECT 141.560000 317.360000 184.760000 318.440000 ;
      RECT 96.560000 317.360000 139.760000 318.440000 ;
      RECT 51.560000 317.360000 94.760000 318.440000 ;
      RECT 6.560000 317.360000 49.760000 318.440000 ;
      RECT 2.530000 317.360000 4.595000 318.440000 ;
      RECT 1.000000 316.490000 199.100000 317.360000 ;
      RECT 0.000000 315.720000 200.100000 316.490000 ;
      RECT 197.570000 315.640000 200.100000 315.720000 ;
      RECT 0.000000 315.640000 2.530000 315.720000 ;
      RECT 197.570000 314.660000 199.100000 315.640000 ;
      RECT 1.000000 314.660000 2.530000 315.640000 ;
      RECT 197.570000 314.640000 200.100000 314.660000 ;
      RECT 188.560000 314.640000 195.770000 315.720000 ;
      RECT 143.560000 314.640000 186.760000 315.720000 ;
      RECT 98.560000 314.640000 141.760000 315.720000 ;
      RECT 53.560000 314.640000 96.760000 315.720000 ;
      RECT 8.560000 314.640000 51.760000 315.720000 ;
      RECT 4.330000 314.640000 6.760000 315.720000 ;
      RECT 0.000000 314.640000 2.530000 314.660000 ;
      RECT 0.000000 314.420000 200.100000 314.640000 ;
      RECT 1.000000 313.440000 199.100000 314.420000 ;
      RECT 0.000000 313.000000 200.100000 313.440000 ;
      RECT 199.370000 312.590000 200.100000 313.000000 ;
      RECT 0.000000 312.590000 0.730000 313.000000 ;
      RECT 186.560000 311.920000 197.570000 313.000000 ;
      RECT 141.560000 311.920000 184.760000 313.000000 ;
      RECT 96.560000 311.920000 139.760000 313.000000 ;
      RECT 51.560000 311.920000 94.760000 313.000000 ;
      RECT 6.560000 311.920000 49.760000 313.000000 ;
      RECT 2.530000 311.920000 4.595000 313.000000 ;
      RECT 1.000000 311.610000 199.100000 311.920000 ;
      RECT 0.000000 311.370000 200.100000 311.610000 ;
      RECT 1.000000 310.390000 199.100000 311.370000 ;
      RECT 0.000000 310.280000 200.100000 310.390000 ;
      RECT 197.570000 309.540000 200.100000 310.280000 ;
      RECT 0.000000 309.540000 2.530000 310.280000 ;
      RECT 197.570000 309.200000 199.100000 309.540000 ;
      RECT 188.560000 309.200000 195.770000 310.280000 ;
      RECT 143.560000 309.200000 186.760000 310.280000 ;
      RECT 98.560000 309.200000 141.760000 310.280000 ;
      RECT 53.560000 309.200000 96.760000 310.280000 ;
      RECT 8.560000 309.200000 51.760000 310.280000 ;
      RECT 4.330000 309.200000 6.760000 310.280000 ;
      RECT 1.000000 309.200000 2.530000 309.540000 ;
      RECT 1.000000 308.560000 199.100000 309.200000 ;
      RECT 0.000000 308.320000 200.100000 308.560000 ;
      RECT 1.000000 307.560000 199.100000 308.320000 ;
      RECT 199.370000 306.490000 200.100000 307.340000 ;
      RECT 0.000000 306.490000 0.730000 307.340000 ;
      RECT 186.560000 306.480000 197.570000 307.560000 ;
      RECT 141.560000 306.480000 184.760000 307.560000 ;
      RECT 96.560000 306.480000 139.760000 307.560000 ;
      RECT 51.560000 306.480000 94.760000 307.560000 ;
      RECT 6.560000 306.480000 49.760000 307.560000 ;
      RECT 2.530000 306.480000 4.595000 307.560000 ;
      RECT 1.000000 305.510000 199.100000 306.480000 ;
      RECT 0.000000 305.270000 200.100000 305.510000 ;
      RECT 1.000000 304.840000 199.100000 305.270000 ;
      RECT 197.570000 304.290000 199.100000 304.840000 ;
      RECT 1.000000 304.290000 2.530000 304.840000 ;
      RECT 197.570000 304.050000 200.100000 304.290000 ;
      RECT 0.000000 304.050000 2.530000 304.290000 ;
      RECT 197.570000 303.760000 199.100000 304.050000 ;
      RECT 188.560000 303.760000 195.770000 304.840000 ;
      RECT 143.560000 303.760000 186.760000 304.840000 ;
      RECT 98.560000 303.760000 141.760000 304.840000 ;
      RECT 53.560000 303.760000 96.760000 304.840000 ;
      RECT 8.560000 303.760000 51.760000 304.840000 ;
      RECT 4.330000 303.760000 6.760000 304.840000 ;
      RECT 1.000000 303.760000 2.530000 304.050000 ;
      RECT 1.000000 303.070000 199.100000 303.760000 ;
      RECT 0.000000 302.220000 200.100000 303.070000 ;
      RECT 1.000000 302.120000 199.100000 302.220000 ;
      RECT 199.370000 301.040000 200.100000 301.240000 ;
      RECT 186.560000 301.040000 197.570000 302.120000 ;
      RECT 141.560000 301.040000 184.760000 302.120000 ;
      RECT 96.560000 301.040000 139.760000 302.120000 ;
      RECT 51.560000 301.040000 94.760000 302.120000 ;
      RECT 6.560000 301.040000 49.760000 302.120000 ;
      RECT 2.530000 301.040000 4.595000 302.120000 ;
      RECT 0.000000 301.040000 0.730000 301.240000 ;
      RECT 0.000000 301.000000 200.100000 301.040000 ;
      RECT 1.000000 300.020000 199.100000 301.000000 ;
      RECT 0.000000 299.400000 200.100000 300.020000 ;
      RECT 197.570000 299.170000 200.100000 299.400000 ;
      RECT 0.000000 299.170000 2.530000 299.400000 ;
      RECT 197.570000 298.320000 199.100000 299.170000 ;
      RECT 188.560000 298.320000 195.770000 299.400000 ;
      RECT 143.560000 298.320000 186.760000 299.400000 ;
      RECT 98.560000 298.320000 141.760000 299.400000 ;
      RECT 53.560000 298.320000 96.760000 299.400000 ;
      RECT 8.560000 298.320000 51.760000 299.400000 ;
      RECT 4.330000 298.320000 6.760000 299.400000 ;
      RECT 1.000000 298.320000 2.530000 299.170000 ;
      RECT 1.000000 298.190000 199.100000 298.320000 ;
      RECT 0.000000 297.950000 200.100000 298.190000 ;
      RECT 1.000000 296.970000 199.100000 297.950000 ;
      RECT 0.000000 296.680000 200.100000 296.970000 ;
      RECT 199.370000 296.120000 200.100000 296.680000 ;
      RECT 0.000000 296.120000 0.730000 296.680000 ;
      RECT 186.560000 295.600000 197.570000 296.680000 ;
      RECT 141.560000 295.600000 184.760000 296.680000 ;
      RECT 96.560000 295.600000 139.760000 296.680000 ;
      RECT 51.560000 295.600000 94.760000 296.680000 ;
      RECT 6.560000 295.600000 49.760000 296.680000 ;
      RECT 2.530000 295.600000 4.595000 296.680000 ;
      RECT 1.000000 295.140000 199.100000 295.600000 ;
      RECT 0.000000 294.900000 200.100000 295.140000 ;
      RECT 1.000000 293.960000 199.100000 294.900000 ;
      RECT 197.570000 293.920000 199.100000 293.960000 ;
      RECT 1.000000 293.920000 2.530000 293.960000 ;
      RECT 197.570000 293.680000 200.100000 293.920000 ;
      RECT 0.000000 293.680000 2.530000 293.920000 ;
      RECT 197.570000 292.880000 199.100000 293.680000 ;
      RECT 188.560000 292.880000 195.770000 293.960000 ;
      RECT 143.560000 292.880000 186.760000 293.960000 ;
      RECT 98.560000 292.880000 141.760000 293.960000 ;
      RECT 53.560000 292.880000 96.760000 293.960000 ;
      RECT 8.560000 292.880000 51.760000 293.960000 ;
      RECT 4.330000 292.880000 6.760000 293.960000 ;
      RECT 1.000000 292.880000 2.530000 293.680000 ;
      RECT 1.000000 292.700000 199.100000 292.880000 ;
      RECT 0.000000 291.850000 200.100000 292.700000 ;
      RECT 1.000000 291.240000 199.100000 291.850000 ;
      RECT 199.370000 290.630000 200.100000 290.870000 ;
      RECT 0.000000 290.630000 0.730000 290.870000 ;
      RECT 186.560000 290.160000 197.570000 291.240000 ;
      RECT 141.560000 290.160000 184.760000 291.240000 ;
      RECT 96.560000 290.160000 139.760000 291.240000 ;
      RECT 51.560000 290.160000 94.760000 291.240000 ;
      RECT 6.560000 290.160000 49.760000 291.240000 ;
      RECT 2.530000 290.160000 4.595000 291.240000 ;
      RECT 1.000000 289.650000 199.100000 290.160000 ;
      RECT 0.000000 288.800000 200.100000 289.650000 ;
      RECT 1.000000 288.520000 199.100000 288.800000 ;
      RECT 197.570000 287.820000 199.100000 288.520000 ;
      RECT 1.000000 287.820000 2.530000 288.520000 ;
      RECT 197.570000 287.580000 200.100000 287.820000 ;
      RECT 0.000000 287.580000 2.530000 287.820000 ;
      RECT 197.570000 287.440000 199.100000 287.580000 ;
      RECT 188.560000 287.440000 195.770000 288.520000 ;
      RECT 143.560000 287.440000 186.760000 288.520000 ;
      RECT 98.560000 287.440000 141.760000 288.520000 ;
      RECT 53.560000 287.440000 96.760000 288.520000 ;
      RECT 8.560000 287.440000 51.760000 288.520000 ;
      RECT 4.330000 287.440000 6.760000 288.520000 ;
      RECT 1.000000 287.440000 2.530000 287.580000 ;
      RECT 1.000000 286.600000 199.100000 287.440000 ;
      RECT 0.000000 285.800000 200.100000 286.600000 ;
      RECT 199.370000 285.750000 200.100000 285.800000 ;
      RECT 0.000000 285.750000 0.730000 285.800000 ;
      RECT 199.370000 284.720000 200.100000 284.770000 ;
      RECT 186.560000 284.720000 197.570000 285.800000 ;
      RECT 141.560000 284.720000 184.760000 285.800000 ;
      RECT 96.560000 284.720000 139.760000 285.800000 ;
      RECT 51.560000 284.720000 94.760000 285.800000 ;
      RECT 6.560000 284.720000 49.760000 285.800000 ;
      RECT 2.530000 284.720000 4.595000 285.800000 ;
      RECT 0.000000 284.720000 0.730000 284.770000 ;
      RECT 0.000000 284.530000 200.100000 284.720000 ;
      RECT 1.000000 283.550000 199.100000 284.530000 ;
      RECT 0.000000 283.080000 200.100000 283.550000 ;
      RECT 197.570000 282.700000 200.100000 283.080000 ;
      RECT 0.000000 282.700000 2.530000 283.080000 ;
      RECT 197.570000 282.000000 199.100000 282.700000 ;
      RECT 188.560000 282.000000 195.770000 283.080000 ;
      RECT 143.560000 282.000000 186.760000 283.080000 ;
      RECT 98.560000 282.000000 141.760000 283.080000 ;
      RECT 53.560000 282.000000 96.760000 283.080000 ;
      RECT 8.560000 282.000000 51.760000 283.080000 ;
      RECT 4.330000 282.000000 6.760000 283.080000 ;
      RECT 1.000000 282.000000 2.530000 282.700000 ;
      RECT 1.000000 281.720000 199.100000 282.000000 ;
      RECT 0.000000 281.480000 200.100000 281.720000 ;
      RECT 1.000000 280.500000 199.100000 281.480000 ;
      RECT 0.000000 280.360000 200.100000 280.500000 ;
      RECT 199.370000 280.260000 200.100000 280.360000 ;
      RECT 0.000000 280.260000 0.730000 280.360000 ;
      RECT 186.560000 279.280000 197.570000 280.360000 ;
      RECT 141.560000 279.280000 184.760000 280.360000 ;
      RECT 96.560000 279.280000 139.760000 280.360000 ;
      RECT 51.560000 279.280000 94.760000 280.360000 ;
      RECT 6.560000 279.280000 49.760000 280.360000 ;
      RECT 2.530000 279.280000 4.595000 280.360000 ;
      RECT 0.000000 278.430000 200.100000 279.280000 ;
      RECT 1.000000 277.640000 199.100000 278.430000 ;
      RECT 197.570000 277.450000 199.100000 277.640000 ;
      RECT 1.000000 277.450000 2.530000 277.640000 ;
      RECT 197.570000 277.210000 200.100000 277.450000 ;
      RECT 0.000000 277.210000 2.530000 277.450000 ;
      RECT 197.570000 276.560000 199.100000 277.210000 ;
      RECT 188.560000 276.560000 195.770000 277.640000 ;
      RECT 143.560000 276.560000 186.760000 277.640000 ;
      RECT 98.560000 276.560000 141.760000 277.640000 ;
      RECT 53.560000 276.560000 96.760000 277.640000 ;
      RECT 8.560000 276.560000 51.760000 277.640000 ;
      RECT 4.330000 276.560000 6.760000 277.640000 ;
      RECT 1.000000 276.560000 2.530000 277.210000 ;
      RECT 1.000000 276.230000 199.100000 276.560000 ;
      RECT 0.000000 275.380000 200.100000 276.230000 ;
      RECT 1.000000 274.920000 199.100000 275.380000 ;
      RECT 199.370000 274.160000 200.100000 274.400000 ;
      RECT 0.000000 274.160000 0.730000 274.400000 ;
      RECT 186.560000 273.840000 197.570000 274.920000 ;
      RECT 141.560000 273.840000 184.760000 274.920000 ;
      RECT 96.560000 273.840000 139.760000 274.920000 ;
      RECT 51.560000 273.840000 94.760000 274.920000 ;
      RECT 6.560000 273.840000 49.760000 274.920000 ;
      RECT 2.530000 273.840000 4.595000 274.920000 ;
      RECT 1.000000 273.180000 199.100000 273.840000 ;
      RECT 0.000000 272.330000 200.100000 273.180000 ;
      RECT 1.000000 272.200000 199.100000 272.330000 ;
      RECT 197.570000 271.350000 199.100000 272.200000 ;
      RECT 1.000000 271.350000 2.530000 272.200000 ;
      RECT 197.570000 271.120000 200.100000 271.350000 ;
      RECT 188.560000 271.120000 195.770000 272.200000 ;
      RECT 143.560000 271.120000 186.760000 272.200000 ;
      RECT 98.560000 271.120000 141.760000 272.200000 ;
      RECT 53.560000 271.120000 96.760000 272.200000 ;
      RECT 8.560000 271.120000 51.760000 272.200000 ;
      RECT 4.330000 271.120000 6.760000 272.200000 ;
      RECT 0.000000 271.120000 2.530000 271.350000 ;
      RECT 0.000000 271.110000 200.100000 271.120000 ;
      RECT 1.000000 270.130000 199.100000 271.110000 ;
      RECT 0.000000 269.480000 200.100000 270.130000 ;
      RECT 199.370000 269.280000 200.100000 269.480000 ;
      RECT 0.000000 269.280000 0.730000 269.480000 ;
      RECT 186.560000 268.400000 197.570000 269.480000 ;
      RECT 141.560000 268.400000 184.760000 269.480000 ;
      RECT 96.560000 268.400000 139.760000 269.480000 ;
      RECT 51.560000 268.400000 94.760000 269.480000 ;
      RECT 6.560000 268.400000 49.760000 269.480000 ;
      RECT 2.530000 268.400000 4.595000 269.480000 ;
      RECT 1.000000 268.300000 199.100000 268.400000 ;
      RECT 0.000000 268.060000 200.100000 268.300000 ;
      RECT 1.000000 267.080000 199.100000 268.060000 ;
      RECT 0.000000 266.840000 200.100000 267.080000 ;
      RECT 1.000000 266.760000 199.100000 266.840000 ;
      RECT 197.570000 265.860000 199.100000 266.760000 ;
      RECT 1.000000 265.860000 2.530000 266.760000 ;
      RECT 197.570000 265.680000 200.100000 265.860000 ;
      RECT 188.560000 265.680000 195.770000 266.760000 ;
      RECT 143.560000 265.680000 186.760000 266.760000 ;
      RECT 98.560000 265.680000 141.760000 266.760000 ;
      RECT 53.560000 265.680000 96.760000 266.760000 ;
      RECT 8.560000 265.680000 51.760000 266.760000 ;
      RECT 4.330000 265.680000 6.760000 266.760000 ;
      RECT 0.000000 265.680000 2.530000 265.860000 ;
      RECT 0.000000 265.010000 200.100000 265.680000 ;
      RECT 1.000000 264.040000 199.100000 265.010000 ;
      RECT 199.370000 263.790000 200.100000 264.030000 ;
      RECT 0.000000 263.790000 0.730000 264.030000 ;
      RECT 186.560000 262.960000 197.570000 264.040000 ;
      RECT 141.560000 262.960000 184.760000 264.040000 ;
      RECT 96.560000 262.960000 139.760000 264.040000 ;
      RECT 51.560000 262.960000 94.760000 264.040000 ;
      RECT 6.560000 262.960000 49.760000 264.040000 ;
      RECT 2.530000 262.960000 4.595000 264.040000 ;
      RECT 1.000000 262.810000 199.100000 262.960000 ;
      RECT 0.000000 261.960000 200.100000 262.810000 ;
      RECT 1.000000 261.320000 199.100000 261.960000 ;
      RECT 197.570000 260.980000 199.100000 261.320000 ;
      RECT 1.000000 260.980000 2.530000 261.320000 ;
      RECT 197.570000 260.740000 200.100000 260.980000 ;
      RECT 0.000000 260.740000 2.530000 260.980000 ;
      RECT 197.570000 260.240000 199.100000 260.740000 ;
      RECT 188.560000 260.240000 195.770000 261.320000 ;
      RECT 143.560000 260.240000 186.760000 261.320000 ;
      RECT 98.560000 260.240000 141.760000 261.320000 ;
      RECT 53.560000 260.240000 96.760000 261.320000 ;
      RECT 8.560000 260.240000 51.760000 261.320000 ;
      RECT 4.330000 260.240000 6.760000 261.320000 ;
      RECT 1.000000 260.240000 2.530000 260.740000 ;
      RECT 1.000000 259.760000 199.100000 260.240000 ;
      RECT 0.000000 258.910000 200.100000 259.760000 ;
      RECT 1.000000 258.600000 199.100000 258.910000 ;
      RECT 199.370000 257.690000 200.100000 257.930000 ;
      RECT 0.000000 257.690000 0.730000 257.930000 ;
      RECT 186.560000 257.520000 197.570000 258.600000 ;
      RECT 141.560000 257.520000 184.760000 258.600000 ;
      RECT 96.560000 257.520000 139.760000 258.600000 ;
      RECT 51.560000 257.520000 94.760000 258.600000 ;
      RECT 6.560000 257.520000 49.760000 258.600000 ;
      RECT 2.530000 257.520000 4.595000 258.600000 ;
      RECT 1.000000 256.710000 199.100000 257.520000 ;
      RECT 0.000000 255.880000 200.100000 256.710000 ;
      RECT 197.570000 255.860000 200.100000 255.880000 ;
      RECT 0.000000 255.860000 2.530000 255.880000 ;
      RECT 197.570000 254.880000 199.100000 255.860000 ;
      RECT 1.000000 254.880000 2.530000 255.860000 ;
      RECT 197.570000 254.800000 200.100000 254.880000 ;
      RECT 188.560000 254.800000 195.770000 255.880000 ;
      RECT 143.560000 254.800000 186.760000 255.880000 ;
      RECT 98.560000 254.800000 141.760000 255.880000 ;
      RECT 53.560000 254.800000 96.760000 255.880000 ;
      RECT 8.560000 254.800000 51.760000 255.880000 ;
      RECT 4.330000 254.800000 6.760000 255.880000 ;
      RECT 0.000000 254.800000 2.530000 254.880000 ;
      RECT 0.000000 254.640000 200.100000 254.800000 ;
      RECT 1.000000 253.660000 199.100000 254.640000 ;
      RECT 0.000000 253.420000 200.100000 253.660000 ;
      RECT 1.000000 253.160000 199.100000 253.420000 ;
      RECT 199.370000 252.080000 200.100000 252.440000 ;
      RECT 186.560000 252.080000 197.570000 253.160000 ;
      RECT 141.560000 252.080000 184.760000 253.160000 ;
      RECT 96.560000 252.080000 139.760000 253.160000 ;
      RECT 51.560000 252.080000 94.760000 253.160000 ;
      RECT 6.560000 252.080000 49.760000 253.160000 ;
      RECT 2.530000 252.080000 4.595000 253.160000 ;
      RECT 0.000000 252.080000 0.730000 252.440000 ;
      RECT 0.000000 251.590000 200.100000 252.080000 ;
      RECT 1.000000 250.610000 199.100000 251.590000 ;
      RECT 0.000000 250.440000 200.100000 250.610000 ;
      RECT 197.570000 250.370000 200.100000 250.440000 ;
      RECT 0.000000 250.370000 2.530000 250.440000 ;
      RECT 197.570000 249.390000 199.100000 250.370000 ;
      RECT 1.000000 249.390000 2.530000 250.370000 ;
      RECT 197.570000 249.360000 200.100000 249.390000 ;
      RECT 188.560000 249.360000 195.770000 250.440000 ;
      RECT 143.560000 249.360000 186.760000 250.440000 ;
      RECT 98.560000 249.360000 141.760000 250.440000 ;
      RECT 53.560000 249.360000 96.760000 250.440000 ;
      RECT 8.560000 249.360000 51.760000 250.440000 ;
      RECT 4.330000 249.360000 6.760000 250.440000 ;
      RECT 0.000000 249.360000 2.530000 249.390000 ;
      RECT 0.000000 248.540000 200.100000 249.360000 ;
      RECT 1.000000 247.720000 199.100000 248.540000 ;
      RECT 199.370000 247.320000 200.100000 247.560000 ;
      RECT 0.000000 247.320000 0.730000 247.560000 ;
      RECT 186.560000 246.640000 197.570000 247.720000 ;
      RECT 141.560000 246.640000 184.760000 247.720000 ;
      RECT 96.560000 246.640000 139.760000 247.720000 ;
      RECT 51.560000 246.640000 94.760000 247.720000 ;
      RECT 6.560000 246.640000 49.760000 247.720000 ;
      RECT 2.530000 246.640000 4.595000 247.720000 ;
      RECT 1.000000 246.340000 199.100000 246.640000 ;
      RECT 0.000000 245.490000 200.100000 246.340000 ;
      RECT 1.000000 245.000000 199.100000 245.490000 ;
      RECT 197.570000 244.510000 199.100000 245.000000 ;
      RECT 1.000000 244.510000 2.530000 245.000000 ;
      RECT 197.570000 244.270000 200.100000 244.510000 ;
      RECT 0.000000 244.270000 2.530000 244.510000 ;
      RECT 197.570000 243.920000 199.100000 244.270000 ;
      RECT 188.560000 243.920000 195.770000 245.000000 ;
      RECT 143.560000 243.920000 186.760000 245.000000 ;
      RECT 98.560000 243.920000 141.760000 245.000000 ;
      RECT 53.560000 243.920000 96.760000 245.000000 ;
      RECT 8.560000 243.920000 51.760000 245.000000 ;
      RECT 4.330000 243.920000 6.760000 245.000000 ;
      RECT 1.000000 243.920000 2.530000 244.270000 ;
      RECT 1.000000 243.290000 199.100000 243.920000 ;
      RECT 0.000000 243.050000 200.100000 243.290000 ;
      RECT 1.000000 242.280000 199.100000 243.050000 ;
      RECT 199.370000 241.220000 200.100000 242.070000 ;
      RECT 0.000000 241.220000 0.730000 242.070000 ;
      RECT 186.560000 241.200000 197.570000 242.280000 ;
      RECT 141.560000 241.200000 184.760000 242.280000 ;
      RECT 96.560000 241.200000 139.760000 242.280000 ;
      RECT 51.560000 241.200000 94.760000 242.280000 ;
      RECT 6.560000 241.200000 49.760000 242.280000 ;
      RECT 2.530000 241.200000 4.595000 242.280000 ;
      RECT 1.000000 240.240000 199.100000 241.200000 ;
      RECT 0.000000 240.000000 200.100000 240.240000 ;
      RECT 1.000000 239.560000 199.100000 240.000000 ;
      RECT 197.570000 239.020000 199.100000 239.560000 ;
      RECT 1.000000 239.020000 2.530000 239.560000 ;
      RECT 197.570000 238.480000 200.100000 239.020000 ;
      RECT 188.560000 238.480000 195.770000 239.560000 ;
      RECT 143.560000 238.480000 186.760000 239.560000 ;
      RECT 98.560000 238.480000 141.760000 239.560000 ;
      RECT 53.560000 238.480000 96.760000 239.560000 ;
      RECT 8.560000 238.480000 51.760000 239.560000 ;
      RECT 4.330000 238.480000 6.760000 239.560000 ;
      RECT 0.000000 238.480000 2.530000 239.020000 ;
      RECT 0.000000 238.170000 200.100000 238.480000 ;
      RECT 1.000000 237.190000 199.100000 238.170000 ;
      RECT 0.000000 236.950000 200.100000 237.190000 ;
      RECT 1.000000 236.840000 199.100000 236.950000 ;
      RECT 199.370000 235.760000 200.100000 235.970000 ;
      RECT 186.560000 235.760000 197.570000 236.840000 ;
      RECT 141.560000 235.760000 184.760000 236.840000 ;
      RECT 96.560000 235.760000 139.760000 236.840000 ;
      RECT 51.560000 235.760000 94.760000 236.840000 ;
      RECT 6.560000 235.760000 49.760000 236.840000 ;
      RECT 2.530000 235.760000 4.595000 236.840000 ;
      RECT 0.000000 235.760000 0.730000 235.970000 ;
      RECT 0.000000 235.120000 200.100000 235.760000 ;
      RECT 1.000000 234.140000 199.100000 235.120000 ;
      RECT 0.000000 234.120000 200.100000 234.140000 ;
      RECT 197.570000 233.900000 200.100000 234.120000 ;
      RECT 0.000000 233.900000 2.530000 234.120000 ;
      RECT 197.570000 233.040000 199.100000 233.900000 ;
      RECT 188.560000 233.040000 195.770000 234.120000 ;
      RECT 143.560000 233.040000 186.760000 234.120000 ;
      RECT 98.560000 233.040000 141.760000 234.120000 ;
      RECT 53.560000 233.040000 96.760000 234.120000 ;
      RECT 8.560000 233.040000 51.760000 234.120000 ;
      RECT 4.330000 233.040000 6.760000 234.120000 ;
      RECT 1.000000 233.040000 2.530000 233.900000 ;
      RECT 1.000000 232.920000 199.100000 233.040000 ;
      RECT 0.000000 232.070000 200.100000 232.920000 ;
      RECT 1.000000 231.400000 199.100000 232.070000 ;
      RECT 199.370000 230.850000 200.100000 231.090000 ;
      RECT 0.000000 230.850000 0.730000 231.090000 ;
      RECT 186.560000 230.320000 197.570000 231.400000 ;
      RECT 141.560000 230.320000 184.760000 231.400000 ;
      RECT 96.560000 230.320000 139.760000 231.400000 ;
      RECT 51.560000 230.320000 94.760000 231.400000 ;
      RECT 6.560000 230.320000 49.760000 231.400000 ;
      RECT 2.530000 230.320000 4.595000 231.400000 ;
      RECT 1.000000 229.870000 199.100000 230.320000 ;
      RECT 0.000000 229.630000 200.100000 229.870000 ;
      RECT 1.000000 228.680000 199.100000 229.630000 ;
      RECT 197.570000 228.650000 199.100000 228.680000 ;
      RECT 1.000000 228.650000 2.530000 228.680000 ;
      RECT 197.570000 227.800000 200.100000 228.650000 ;
      RECT 0.000000 227.800000 2.530000 228.650000 ;
      RECT 197.570000 227.600000 199.100000 227.800000 ;
      RECT 188.560000 227.600000 195.770000 228.680000 ;
      RECT 143.560000 227.600000 186.760000 228.680000 ;
      RECT 98.560000 227.600000 141.760000 228.680000 ;
      RECT 53.560000 227.600000 96.760000 228.680000 ;
      RECT 8.560000 227.600000 51.760000 228.680000 ;
      RECT 4.330000 227.600000 6.760000 228.680000 ;
      RECT 1.000000 227.600000 2.530000 227.800000 ;
      RECT 1.000000 226.820000 199.100000 227.600000 ;
      RECT 0.000000 226.580000 200.100000 226.820000 ;
      RECT 1.000000 225.960000 199.100000 226.580000 ;
      RECT 199.370000 224.880000 200.100000 225.600000 ;
      RECT 186.560000 224.880000 197.570000 225.960000 ;
      RECT 141.560000 224.880000 184.760000 225.960000 ;
      RECT 96.560000 224.880000 139.760000 225.960000 ;
      RECT 51.560000 224.880000 94.760000 225.960000 ;
      RECT 6.560000 224.880000 49.760000 225.960000 ;
      RECT 2.530000 224.880000 4.595000 225.960000 ;
      RECT 0.000000 224.880000 0.730000 225.600000 ;
      RECT 0.000000 224.750000 200.100000 224.880000 ;
      RECT 1.000000 223.770000 199.100000 224.750000 ;
      RECT 0.000000 223.530000 200.100000 223.770000 ;
      RECT 1.000000 223.240000 199.100000 223.530000 ;
      RECT 197.570000 222.550000 199.100000 223.240000 ;
      RECT 1.000000 222.550000 2.530000 223.240000 ;
      RECT 197.570000 222.160000 200.100000 222.550000 ;
      RECT 188.560000 222.160000 195.770000 223.240000 ;
      RECT 143.560000 222.160000 186.760000 223.240000 ;
      RECT 98.560000 222.160000 141.760000 223.240000 ;
      RECT 53.560000 222.160000 96.760000 223.240000 ;
      RECT 8.560000 222.160000 51.760000 223.240000 ;
      RECT 4.330000 222.160000 6.760000 223.240000 ;
      RECT 0.000000 222.160000 2.530000 222.550000 ;
      RECT 0.000000 221.700000 200.100000 222.160000 ;
      RECT 1.000000 220.720000 199.100000 221.700000 ;
      RECT 0.000000 220.520000 200.100000 220.720000 ;
      RECT 199.370000 220.480000 200.100000 220.520000 ;
      RECT 0.000000 220.480000 0.730000 220.520000 ;
      RECT 199.370000 219.440000 200.100000 219.500000 ;
      RECT 186.560000 219.440000 197.570000 220.520000 ;
      RECT 141.560000 219.440000 184.760000 220.520000 ;
      RECT 96.560000 219.440000 139.760000 220.520000 ;
      RECT 51.560000 219.440000 94.760000 220.520000 ;
      RECT 6.560000 219.440000 49.760000 220.520000 ;
      RECT 2.530000 219.440000 4.595000 220.520000 ;
      RECT 0.000000 219.440000 0.730000 219.500000 ;
      RECT 0.000000 218.650000 200.100000 219.440000 ;
      RECT 1.000000 217.800000 199.100000 218.650000 ;
      RECT 197.570000 217.670000 199.100000 217.800000 ;
      RECT 1.000000 217.670000 2.530000 217.800000 ;
      RECT 197.570000 217.430000 200.100000 217.670000 ;
      RECT 0.000000 217.430000 2.530000 217.670000 ;
      RECT 197.570000 216.720000 199.100000 217.430000 ;
      RECT 188.560000 216.720000 195.770000 217.800000 ;
      RECT 143.560000 216.720000 186.760000 217.800000 ;
      RECT 98.560000 216.720000 141.760000 217.800000 ;
      RECT 53.560000 216.720000 96.760000 217.800000 ;
      RECT 8.560000 216.720000 51.760000 217.800000 ;
      RECT 4.330000 216.720000 6.760000 217.800000 ;
      RECT 1.000000 216.720000 2.530000 217.430000 ;
      RECT 1.000000 216.450000 199.100000 216.720000 ;
      RECT 0.000000 216.210000 200.100000 216.450000 ;
      RECT 1.000000 215.230000 199.100000 216.210000 ;
      RECT 0.000000 215.080000 200.100000 215.230000 ;
      RECT 199.370000 214.380000 200.100000 215.080000 ;
      RECT 0.000000 214.380000 0.730000 215.080000 ;
      RECT 186.560000 214.000000 197.570000 215.080000 ;
      RECT 141.560000 214.000000 184.760000 215.080000 ;
      RECT 96.560000 214.000000 139.760000 215.080000 ;
      RECT 51.560000 214.000000 94.760000 215.080000 ;
      RECT 6.560000 214.000000 49.760000 215.080000 ;
      RECT 2.530000 214.000000 4.595000 215.080000 ;
      RECT 1.000000 213.400000 199.100000 214.000000 ;
      RECT 0.000000 213.160000 200.100000 213.400000 ;
      RECT 1.000000 212.360000 199.100000 213.160000 ;
      RECT 197.570000 212.180000 199.100000 212.360000 ;
      RECT 1.000000 212.180000 2.530000 212.360000 ;
      RECT 197.570000 211.330000 200.100000 212.180000 ;
      RECT 0.000000 211.330000 2.530000 212.180000 ;
      RECT 197.570000 211.280000 199.100000 211.330000 ;
      RECT 188.560000 211.280000 195.770000 212.360000 ;
      RECT 143.560000 211.280000 186.760000 212.360000 ;
      RECT 98.560000 211.280000 141.760000 212.360000 ;
      RECT 53.560000 211.280000 96.760000 212.360000 ;
      RECT 8.560000 211.280000 51.760000 212.360000 ;
      RECT 4.330000 211.280000 6.760000 212.360000 ;
      RECT 1.000000 211.280000 2.530000 211.330000 ;
      RECT 1.000000 210.350000 199.100000 211.280000 ;
      RECT 0.000000 210.110000 200.100000 210.350000 ;
      RECT 1.000000 209.640000 199.100000 210.110000 ;
      RECT 199.370000 208.560000 200.100000 209.130000 ;
      RECT 186.560000 208.560000 197.570000 209.640000 ;
      RECT 141.560000 208.560000 184.760000 209.640000 ;
      RECT 96.560000 208.560000 139.760000 209.640000 ;
      RECT 51.560000 208.560000 94.760000 209.640000 ;
      RECT 6.560000 208.560000 49.760000 209.640000 ;
      RECT 2.530000 208.560000 4.595000 209.640000 ;
      RECT 0.000000 208.560000 0.730000 209.130000 ;
      RECT 0.000000 208.280000 200.100000 208.560000 ;
      RECT 1.000000 207.300000 199.100000 208.280000 ;
      RECT 0.000000 207.060000 200.100000 207.300000 ;
      RECT 1.000000 206.920000 199.100000 207.060000 ;
      RECT 197.570000 206.080000 199.100000 206.920000 ;
      RECT 1.000000 206.080000 2.530000 206.920000 ;
      RECT 197.570000 205.840000 200.100000 206.080000 ;
      RECT 188.560000 205.840000 195.770000 206.920000 ;
      RECT 143.560000 205.840000 186.760000 206.920000 ;
      RECT 98.560000 205.840000 141.760000 206.920000 ;
      RECT 53.560000 205.840000 96.760000 206.920000 ;
      RECT 8.560000 205.840000 51.760000 206.920000 ;
      RECT 4.330000 205.840000 6.760000 206.920000 ;
      RECT 0.000000 205.840000 2.530000 206.080000 ;
      RECT 1.000000 204.860000 199.100000 205.840000 ;
      RECT 0.000000 204.200000 200.100000 204.860000 ;
      RECT 199.370000 203.120000 200.100000 204.200000 ;
      RECT 186.560000 203.120000 197.570000 204.200000 ;
      RECT 141.560000 203.120000 184.760000 204.200000 ;
      RECT 96.560000 203.120000 139.760000 204.200000 ;
      RECT 51.560000 203.120000 94.760000 204.200000 ;
      RECT 6.560000 203.120000 49.760000 204.200000 ;
      RECT 2.530000 203.120000 4.595000 204.200000 ;
      RECT 0.000000 203.120000 0.730000 204.200000 ;
      RECT 0.000000 201.480000 200.100000 203.120000 ;
      RECT 197.570000 200.400000 200.100000 201.480000 ;
      RECT 188.560000 200.400000 195.770000 201.480000 ;
      RECT 143.560000 200.400000 186.760000 201.480000 ;
      RECT 98.560000 200.400000 141.760000 201.480000 ;
      RECT 53.560000 200.400000 96.760000 201.480000 ;
      RECT 8.560000 200.400000 51.760000 201.480000 ;
      RECT 4.330000 200.400000 6.760000 201.480000 ;
      RECT 0.000000 200.400000 2.530000 201.480000 ;
      RECT 0.000000 198.760000 200.100000 200.400000 ;
      RECT 199.370000 197.680000 200.100000 198.760000 ;
      RECT 186.560000 197.680000 197.570000 198.760000 ;
      RECT 141.560000 197.680000 184.760000 198.760000 ;
      RECT 96.560000 197.680000 139.760000 198.760000 ;
      RECT 51.560000 197.680000 94.760000 198.760000 ;
      RECT 6.560000 197.680000 49.760000 198.760000 ;
      RECT 2.530000 197.680000 4.595000 198.760000 ;
      RECT 0.000000 197.680000 0.730000 198.760000 ;
      RECT 0.000000 196.040000 200.100000 197.680000 ;
      RECT 197.570000 195.470000 200.100000 196.040000 ;
      RECT 0.000000 195.470000 2.530000 196.040000 ;
      RECT 197.570000 194.960000 199.100000 195.470000 ;
      RECT 188.560000 194.960000 195.770000 196.040000 ;
      RECT 143.560000 194.960000 186.760000 196.040000 ;
      RECT 98.560000 194.960000 141.760000 196.040000 ;
      RECT 53.560000 194.960000 96.760000 196.040000 ;
      RECT 8.560000 194.960000 51.760000 196.040000 ;
      RECT 4.330000 194.960000 6.760000 196.040000 ;
      RECT 1.000000 194.960000 2.530000 195.470000 ;
      RECT 1.000000 194.490000 199.100000 194.960000 ;
      RECT 0.000000 193.640000 200.100000 194.490000 ;
      RECT 1.000000 193.320000 199.100000 193.640000 ;
      RECT 199.370000 192.420000 200.100000 192.660000 ;
      RECT 0.000000 192.420000 0.730000 192.660000 ;
      RECT 186.560000 192.240000 197.570000 193.320000 ;
      RECT 141.560000 192.240000 184.760000 193.320000 ;
      RECT 96.560000 192.240000 139.760000 193.320000 ;
      RECT 51.560000 192.240000 94.760000 193.320000 ;
      RECT 6.560000 192.240000 49.760000 193.320000 ;
      RECT 2.530000 192.240000 4.595000 193.320000 ;
      RECT 1.000000 191.440000 199.100000 192.240000 ;
      RECT 0.000000 190.600000 200.100000 191.440000 ;
      RECT 197.570000 190.590000 200.100000 190.600000 ;
      RECT 0.000000 190.590000 2.530000 190.600000 ;
      RECT 197.570000 189.610000 199.100000 190.590000 ;
      RECT 1.000000 189.610000 2.530000 190.590000 ;
      RECT 197.570000 189.520000 200.100000 189.610000 ;
      RECT 188.560000 189.520000 195.770000 190.600000 ;
      RECT 143.560000 189.520000 186.760000 190.600000 ;
      RECT 98.560000 189.520000 141.760000 190.600000 ;
      RECT 53.560000 189.520000 96.760000 190.600000 ;
      RECT 8.560000 189.520000 51.760000 190.600000 ;
      RECT 4.330000 189.520000 6.760000 190.600000 ;
      RECT 0.000000 189.520000 2.530000 189.610000 ;
      RECT 0.000000 189.370000 200.100000 189.520000 ;
      RECT 1.000000 188.390000 199.100000 189.370000 ;
      RECT 0.000000 187.880000 200.100000 188.390000 ;
      RECT 199.370000 187.540000 200.100000 187.880000 ;
      RECT 0.000000 187.540000 0.730000 187.880000 ;
      RECT 186.560000 186.800000 197.570000 187.880000 ;
      RECT 141.560000 186.800000 184.760000 187.880000 ;
      RECT 96.560000 186.800000 139.760000 187.880000 ;
      RECT 51.560000 186.800000 94.760000 187.880000 ;
      RECT 6.560000 186.800000 49.760000 187.880000 ;
      RECT 2.530000 186.800000 4.595000 187.880000 ;
      RECT 1.000000 186.560000 199.100000 186.800000 ;
      RECT 0.000000 186.320000 200.100000 186.560000 ;
      RECT 1.000000 185.340000 199.100000 186.320000 ;
      RECT 0.000000 185.160000 200.100000 185.340000 ;
      RECT 197.570000 184.490000 200.100000 185.160000 ;
      RECT 0.000000 184.490000 2.530000 185.160000 ;
      RECT 197.570000 184.080000 199.100000 184.490000 ;
      RECT 188.560000 184.080000 195.770000 185.160000 ;
      RECT 143.560000 184.080000 186.760000 185.160000 ;
      RECT 98.560000 184.080000 141.760000 185.160000 ;
      RECT 53.560000 184.080000 96.760000 185.160000 ;
      RECT 8.560000 184.080000 51.760000 185.160000 ;
      RECT 4.330000 184.080000 6.760000 185.160000 ;
      RECT 1.000000 184.080000 2.530000 184.490000 ;
      RECT 1.000000 183.510000 199.100000 184.080000 ;
      RECT 0.000000 183.270000 200.100000 183.510000 ;
      RECT 1.000000 182.440000 199.100000 183.270000 ;
      RECT 199.370000 181.440000 200.100000 182.290000 ;
      RECT 0.000000 181.440000 0.730000 182.290000 ;
      RECT 186.560000 181.360000 197.570000 182.440000 ;
      RECT 141.560000 181.360000 184.760000 182.440000 ;
      RECT 96.560000 181.360000 139.760000 182.440000 ;
      RECT 51.560000 181.360000 94.760000 182.440000 ;
      RECT 6.560000 181.360000 49.760000 182.440000 ;
      RECT 2.530000 181.360000 4.595000 182.440000 ;
      RECT 1.000000 180.460000 199.100000 181.360000 ;
      RECT 0.000000 180.220000 200.100000 180.460000 ;
      RECT 1.000000 179.720000 199.100000 180.220000 ;
      RECT 197.570000 179.240000 199.100000 179.720000 ;
      RECT 1.000000 179.240000 2.530000 179.720000 ;
      RECT 197.570000 179.000000 200.100000 179.240000 ;
      RECT 0.000000 179.000000 2.530000 179.240000 ;
      RECT 197.570000 178.640000 199.100000 179.000000 ;
      RECT 188.560000 178.640000 195.770000 179.720000 ;
      RECT 143.560000 178.640000 186.760000 179.720000 ;
      RECT 98.560000 178.640000 141.760000 179.720000 ;
      RECT 53.560000 178.640000 96.760000 179.720000 ;
      RECT 8.560000 178.640000 51.760000 179.720000 ;
      RECT 4.330000 178.640000 6.760000 179.720000 ;
      RECT 1.000000 178.640000 2.530000 179.000000 ;
      RECT 1.000000 178.020000 199.100000 178.640000 ;
      RECT 0.000000 177.170000 200.100000 178.020000 ;
      RECT 1.000000 177.000000 199.100000 177.170000 ;
      RECT 199.370000 175.950000 200.100000 176.190000 ;
      RECT 0.000000 175.950000 0.730000 176.190000 ;
      RECT 186.560000 175.920000 197.570000 177.000000 ;
      RECT 141.560000 175.920000 184.760000 177.000000 ;
      RECT 96.560000 175.920000 139.760000 177.000000 ;
      RECT 51.560000 175.920000 94.760000 177.000000 ;
      RECT 6.560000 175.920000 49.760000 177.000000 ;
      RECT 2.530000 175.920000 4.595000 177.000000 ;
      RECT 1.000000 174.970000 199.100000 175.920000 ;
      RECT 0.000000 174.280000 200.100000 174.970000 ;
      RECT 197.570000 174.120000 200.100000 174.280000 ;
      RECT 0.000000 174.120000 2.530000 174.280000 ;
      RECT 197.570000 173.200000 199.100000 174.120000 ;
      RECT 188.560000 173.200000 195.770000 174.280000 ;
      RECT 143.560000 173.200000 186.760000 174.280000 ;
      RECT 98.560000 173.200000 141.760000 174.280000 ;
      RECT 53.560000 173.200000 96.760000 174.280000 ;
      RECT 8.560000 173.200000 51.760000 174.280000 ;
      RECT 4.330000 173.200000 6.760000 174.280000 ;
      RECT 1.000000 173.200000 2.530000 174.120000 ;
      RECT 1.000000 173.140000 199.100000 173.200000 ;
      RECT 0.000000 172.900000 200.100000 173.140000 ;
      RECT 1.000000 171.920000 199.100000 172.900000 ;
      RECT 0.000000 171.560000 200.100000 171.920000 ;
      RECT 199.370000 171.070000 200.100000 171.560000 ;
      RECT 0.000000 171.070000 0.730000 171.560000 ;
      RECT 186.560000 170.480000 197.570000 171.560000 ;
      RECT 141.560000 170.480000 184.760000 171.560000 ;
      RECT 96.560000 170.480000 139.760000 171.560000 ;
      RECT 51.560000 170.480000 94.760000 171.560000 ;
      RECT 6.560000 170.480000 49.760000 171.560000 ;
      RECT 2.530000 170.480000 4.595000 171.560000 ;
      RECT 1.000000 170.090000 199.100000 170.480000 ;
      RECT 0.000000 169.850000 200.100000 170.090000 ;
      RECT 1.000000 168.870000 199.100000 169.850000 ;
      RECT 0.000000 168.840000 200.100000 168.870000 ;
      RECT 197.570000 168.020000 200.100000 168.840000 ;
      RECT 0.000000 168.020000 2.530000 168.840000 ;
      RECT 197.570000 167.760000 199.100000 168.020000 ;
      RECT 188.560000 167.760000 195.770000 168.840000 ;
      RECT 143.560000 167.760000 186.760000 168.840000 ;
      RECT 98.560000 167.760000 141.760000 168.840000 ;
      RECT 53.560000 167.760000 96.760000 168.840000 ;
      RECT 8.560000 167.760000 51.760000 168.840000 ;
      RECT 4.330000 167.760000 6.760000 168.840000 ;
      RECT 1.000000 167.760000 2.530000 168.020000 ;
      RECT 1.000000 167.040000 199.100000 167.760000 ;
      RECT 0.000000 166.800000 200.100000 167.040000 ;
      RECT 1.000000 166.120000 199.100000 166.800000 ;
      RECT 199.370000 165.580000 200.100000 165.820000 ;
      RECT 0.000000 165.580000 0.730000 165.820000 ;
      RECT 186.560000 165.040000 197.570000 166.120000 ;
      RECT 141.560000 165.040000 184.760000 166.120000 ;
      RECT 96.560000 165.040000 139.760000 166.120000 ;
      RECT 51.560000 165.040000 94.760000 166.120000 ;
      RECT 6.560000 165.040000 49.760000 166.120000 ;
      RECT 2.530000 165.040000 4.595000 166.120000 ;
      RECT 1.000000 164.600000 199.100000 165.040000 ;
      RECT 0.000000 163.750000 200.100000 164.600000 ;
      RECT 1.000000 163.400000 199.100000 163.750000 ;
      RECT 197.570000 162.770000 199.100000 163.400000 ;
      RECT 1.000000 162.770000 2.530000 163.400000 ;
      RECT 197.570000 162.530000 200.100000 162.770000 ;
      RECT 0.000000 162.530000 2.530000 162.770000 ;
      RECT 197.570000 162.320000 199.100000 162.530000 ;
      RECT 188.560000 162.320000 195.770000 163.400000 ;
      RECT 143.560000 162.320000 186.760000 163.400000 ;
      RECT 98.560000 162.320000 141.760000 163.400000 ;
      RECT 53.560000 162.320000 96.760000 163.400000 ;
      RECT 8.560000 162.320000 51.760000 163.400000 ;
      RECT 4.330000 162.320000 6.760000 163.400000 ;
      RECT 1.000000 162.320000 2.530000 162.530000 ;
      RECT 1.000000 161.550000 199.100000 162.320000 ;
      RECT 0.000000 160.700000 200.100000 161.550000 ;
      RECT 1.000000 160.680000 199.100000 160.700000 ;
      RECT 199.370000 159.600000 200.100000 159.720000 ;
      RECT 186.560000 159.600000 197.570000 160.680000 ;
      RECT 141.560000 159.600000 184.760000 160.680000 ;
      RECT 96.560000 159.600000 139.760000 160.680000 ;
      RECT 51.560000 159.600000 94.760000 160.680000 ;
      RECT 6.560000 159.600000 49.760000 160.680000 ;
      RECT 2.530000 159.600000 4.595000 160.680000 ;
      RECT 0.000000 159.600000 0.730000 159.720000 ;
      RECT 0.000000 159.480000 200.100000 159.600000 ;
      RECT 1.000000 158.500000 199.100000 159.480000 ;
      RECT 0.000000 157.960000 200.100000 158.500000 ;
      RECT 197.570000 157.650000 200.100000 157.960000 ;
      RECT 0.000000 157.650000 2.530000 157.960000 ;
      RECT 197.570000 156.880000 199.100000 157.650000 ;
      RECT 188.560000 156.880000 195.770000 157.960000 ;
      RECT 143.560000 156.880000 186.760000 157.960000 ;
      RECT 98.560000 156.880000 141.760000 157.960000 ;
      RECT 53.560000 156.880000 96.760000 157.960000 ;
      RECT 8.560000 156.880000 51.760000 157.960000 ;
      RECT 4.330000 156.880000 6.760000 157.960000 ;
      RECT 1.000000 156.880000 2.530000 157.650000 ;
      RECT 1.000000 156.670000 199.100000 156.880000 ;
      RECT 0.000000 156.430000 200.100000 156.670000 ;
      RECT 1.000000 155.450000 199.100000 156.430000 ;
      RECT 0.000000 155.240000 200.100000 155.450000 ;
      RECT 199.370000 154.600000 200.100000 155.240000 ;
      RECT 0.000000 154.600000 0.730000 155.240000 ;
      RECT 186.560000 154.160000 197.570000 155.240000 ;
      RECT 141.560000 154.160000 184.760000 155.240000 ;
      RECT 96.560000 154.160000 139.760000 155.240000 ;
      RECT 51.560000 154.160000 94.760000 155.240000 ;
      RECT 6.560000 154.160000 49.760000 155.240000 ;
      RECT 2.530000 154.160000 4.595000 155.240000 ;
      RECT 1.000000 153.620000 199.100000 154.160000 ;
      RECT 0.000000 153.380000 200.100000 153.620000 ;
      RECT 1.000000 152.520000 199.100000 153.380000 ;
      RECT 197.570000 152.400000 199.100000 152.520000 ;
      RECT 1.000000 152.400000 2.530000 152.520000 ;
      RECT 197.570000 151.550000 200.100000 152.400000 ;
      RECT 0.000000 151.550000 2.530000 152.400000 ;
      RECT 197.570000 151.440000 199.100000 151.550000 ;
      RECT 188.560000 151.440000 195.770000 152.520000 ;
      RECT 143.560000 151.440000 186.760000 152.520000 ;
      RECT 98.560000 151.440000 141.760000 152.520000 ;
      RECT 53.560000 151.440000 96.760000 152.520000 ;
      RECT 8.560000 151.440000 51.760000 152.520000 ;
      RECT 4.330000 151.440000 6.760000 152.520000 ;
      RECT 1.000000 151.440000 2.530000 151.550000 ;
      RECT 1.000000 150.570000 199.100000 151.440000 ;
      RECT 0.000000 150.330000 200.100000 150.570000 ;
      RECT 1.000000 149.800000 199.100000 150.330000 ;
      RECT 199.370000 149.110000 200.100000 149.350000 ;
      RECT 0.000000 149.110000 0.730000 149.350000 ;
      RECT 186.560000 148.720000 197.570000 149.800000 ;
      RECT 141.560000 148.720000 184.760000 149.800000 ;
      RECT 96.560000 148.720000 139.760000 149.800000 ;
      RECT 51.560000 148.720000 94.760000 149.800000 ;
      RECT 6.560000 148.720000 49.760000 149.800000 ;
      RECT 2.530000 148.720000 4.595000 149.800000 ;
      RECT 1.000000 148.130000 199.100000 148.720000 ;
      RECT 0.000000 147.280000 200.100000 148.130000 ;
      RECT 1.000000 147.080000 199.100000 147.280000 ;
      RECT 197.570000 146.300000 199.100000 147.080000 ;
      RECT 1.000000 146.300000 2.530000 147.080000 ;
      RECT 197.570000 146.060000 200.100000 146.300000 ;
      RECT 0.000000 146.060000 2.530000 146.300000 ;
      RECT 197.570000 146.000000 199.100000 146.060000 ;
      RECT 188.560000 146.000000 195.770000 147.080000 ;
      RECT 143.560000 146.000000 186.760000 147.080000 ;
      RECT 98.560000 146.000000 141.760000 147.080000 ;
      RECT 53.560000 146.000000 96.760000 147.080000 ;
      RECT 8.560000 146.000000 51.760000 147.080000 ;
      RECT 4.330000 146.000000 6.760000 147.080000 ;
      RECT 1.000000 146.000000 2.530000 146.060000 ;
      RECT 1.000000 145.080000 199.100000 146.000000 ;
      RECT 0.000000 144.360000 200.100000 145.080000 ;
      RECT 199.370000 144.230000 200.100000 144.360000 ;
      RECT 0.000000 144.230000 0.730000 144.360000 ;
      RECT 186.560000 143.280000 197.570000 144.360000 ;
      RECT 141.560000 143.280000 184.760000 144.360000 ;
      RECT 96.560000 143.280000 139.760000 144.360000 ;
      RECT 51.560000 143.280000 94.760000 144.360000 ;
      RECT 6.560000 143.280000 49.760000 144.360000 ;
      RECT 2.530000 143.280000 4.595000 144.360000 ;
      RECT 1.000000 143.250000 199.100000 143.280000 ;
      RECT 0.000000 143.010000 200.100000 143.250000 ;
      RECT 1.000000 142.030000 199.100000 143.010000 ;
      RECT 0.000000 141.640000 200.100000 142.030000 ;
      RECT 197.570000 141.180000 200.100000 141.640000 ;
      RECT 0.000000 141.180000 2.530000 141.640000 ;
      RECT 197.570000 140.560000 199.100000 141.180000 ;
      RECT 188.560000 140.560000 195.770000 141.640000 ;
      RECT 143.560000 140.560000 186.760000 141.640000 ;
      RECT 98.560000 140.560000 141.760000 141.640000 ;
      RECT 53.560000 140.560000 96.760000 141.640000 ;
      RECT 8.560000 140.560000 51.760000 141.640000 ;
      RECT 4.330000 140.560000 6.760000 141.640000 ;
      RECT 1.000000 140.560000 2.530000 141.180000 ;
      RECT 1.000000 140.200000 199.100000 140.560000 ;
      RECT 0.000000 139.960000 200.100000 140.200000 ;
      RECT 1.000000 138.980000 199.100000 139.960000 ;
      RECT 0.000000 138.920000 200.100000 138.980000 ;
      RECT 199.370000 138.130000 200.100000 138.920000 ;
      RECT 0.000000 138.130000 0.730000 138.920000 ;
      RECT 186.560000 137.840000 197.570000 138.920000 ;
      RECT 141.560000 137.840000 184.760000 138.920000 ;
      RECT 96.560000 137.840000 139.760000 138.920000 ;
      RECT 51.560000 137.840000 94.760000 138.920000 ;
      RECT 6.560000 137.840000 49.760000 138.920000 ;
      RECT 2.530000 137.840000 4.595000 138.920000 ;
      RECT 1.000000 137.150000 199.100000 137.840000 ;
      RECT 0.000000 136.910000 200.100000 137.150000 ;
      RECT 1.000000 136.200000 199.100000 136.910000 ;
      RECT 197.570000 135.930000 199.100000 136.200000 ;
      RECT 1.000000 135.930000 2.530000 136.200000 ;
      RECT 197.570000 135.690000 200.100000 135.930000 ;
      RECT 0.000000 135.690000 2.530000 135.930000 ;
      RECT 197.570000 135.120000 199.100000 135.690000 ;
      RECT 188.560000 135.120000 195.770000 136.200000 ;
      RECT 143.560000 135.120000 186.760000 136.200000 ;
      RECT 98.560000 135.120000 141.760000 136.200000 ;
      RECT 53.560000 135.120000 96.760000 136.200000 ;
      RECT 8.560000 135.120000 51.760000 136.200000 ;
      RECT 4.330000 135.120000 6.760000 136.200000 ;
      RECT 1.000000 135.120000 2.530000 135.690000 ;
      RECT 1.000000 134.710000 199.100000 135.120000 ;
      RECT 0.000000 133.860000 200.100000 134.710000 ;
      RECT 1.000000 133.480000 199.100000 133.860000 ;
      RECT 199.370000 132.640000 200.100000 132.880000 ;
      RECT 0.000000 132.640000 0.730000 132.880000 ;
      RECT 186.560000 132.400000 197.570000 133.480000 ;
      RECT 141.560000 132.400000 184.760000 133.480000 ;
      RECT 96.560000 132.400000 139.760000 133.480000 ;
      RECT 51.560000 132.400000 94.760000 133.480000 ;
      RECT 6.560000 132.400000 49.760000 133.480000 ;
      RECT 2.530000 132.400000 4.595000 133.480000 ;
      RECT 1.000000 131.660000 199.100000 132.400000 ;
      RECT 0.000000 130.810000 200.100000 131.660000 ;
      RECT 1.000000 130.760000 199.100000 130.810000 ;
      RECT 197.570000 129.830000 199.100000 130.760000 ;
      RECT 1.000000 129.830000 2.530000 130.760000 ;
      RECT 197.570000 129.680000 200.100000 129.830000 ;
      RECT 188.560000 129.680000 195.770000 130.760000 ;
      RECT 143.560000 129.680000 186.760000 130.760000 ;
      RECT 98.560000 129.680000 141.760000 130.760000 ;
      RECT 53.560000 129.680000 96.760000 130.760000 ;
      RECT 8.560000 129.680000 51.760000 130.760000 ;
      RECT 4.330000 129.680000 6.760000 130.760000 ;
      RECT 0.000000 129.680000 2.530000 129.830000 ;
      RECT 0.000000 129.590000 200.100000 129.680000 ;
      RECT 1.000000 128.610000 199.100000 129.590000 ;
      RECT 0.000000 128.040000 200.100000 128.610000 ;
      RECT 199.370000 127.760000 200.100000 128.040000 ;
      RECT 0.000000 127.760000 0.730000 128.040000 ;
      RECT 186.560000 126.960000 197.570000 128.040000 ;
      RECT 141.560000 126.960000 184.760000 128.040000 ;
      RECT 96.560000 126.960000 139.760000 128.040000 ;
      RECT 51.560000 126.960000 94.760000 128.040000 ;
      RECT 6.560000 126.960000 49.760000 128.040000 ;
      RECT 2.530000 126.960000 4.595000 128.040000 ;
      RECT 1.000000 126.780000 199.100000 126.960000 ;
      RECT 0.000000 126.540000 200.100000 126.780000 ;
      RECT 1.000000 125.560000 199.100000 126.540000 ;
      RECT 0.000000 125.320000 200.100000 125.560000 ;
      RECT 197.570000 124.710000 200.100000 125.320000 ;
      RECT 0.000000 124.710000 2.530000 125.320000 ;
      RECT 197.570000 124.240000 199.100000 124.710000 ;
      RECT 188.560000 124.240000 195.770000 125.320000 ;
      RECT 143.560000 124.240000 186.760000 125.320000 ;
      RECT 98.560000 124.240000 141.760000 125.320000 ;
      RECT 53.560000 124.240000 96.760000 125.320000 ;
      RECT 8.560000 124.240000 51.760000 125.320000 ;
      RECT 4.330000 124.240000 6.760000 125.320000 ;
      RECT 1.000000 124.240000 2.530000 124.710000 ;
      RECT 1.000000 123.730000 199.100000 124.240000 ;
      RECT 0.000000 123.490000 200.100000 123.730000 ;
      RECT 1.000000 122.600000 199.100000 123.490000 ;
      RECT 199.370000 122.270000 200.100000 122.510000 ;
      RECT 0.000000 122.270000 0.730000 122.510000 ;
      RECT 186.560000 121.520000 197.570000 122.600000 ;
      RECT 141.560000 121.520000 184.760000 122.600000 ;
      RECT 96.560000 121.520000 139.760000 122.600000 ;
      RECT 51.560000 121.520000 94.760000 122.600000 ;
      RECT 6.560000 121.520000 49.760000 122.600000 ;
      RECT 2.530000 121.520000 4.595000 122.600000 ;
      RECT 1.000000 121.290000 199.100000 121.520000 ;
      RECT 0.000000 120.440000 200.100000 121.290000 ;
      RECT 1.000000 119.880000 199.100000 120.440000 ;
      RECT 197.570000 119.460000 199.100000 119.880000 ;
      RECT 1.000000 119.460000 2.530000 119.880000 ;
      RECT 197.570000 119.220000 200.100000 119.460000 ;
      RECT 0.000000 119.220000 2.530000 119.460000 ;
      RECT 197.570000 118.800000 199.100000 119.220000 ;
      RECT 188.560000 118.800000 195.770000 119.880000 ;
      RECT 143.560000 118.800000 186.760000 119.880000 ;
      RECT 98.560000 118.800000 141.760000 119.880000 ;
      RECT 53.560000 118.800000 96.760000 119.880000 ;
      RECT 8.560000 118.800000 51.760000 119.880000 ;
      RECT 4.330000 118.800000 6.760000 119.880000 ;
      RECT 1.000000 118.800000 2.530000 119.220000 ;
      RECT 1.000000 118.240000 199.100000 118.800000 ;
      RECT 0.000000 117.390000 200.100000 118.240000 ;
      RECT 1.000000 117.160000 199.100000 117.390000 ;
      RECT 199.370000 116.170000 200.100000 116.410000 ;
      RECT 0.000000 116.170000 0.730000 116.410000 ;
      RECT 186.560000 116.080000 197.570000 117.160000 ;
      RECT 141.560000 116.080000 184.760000 117.160000 ;
      RECT 96.560000 116.080000 139.760000 117.160000 ;
      RECT 51.560000 116.080000 94.760000 117.160000 ;
      RECT 6.560000 116.080000 49.760000 117.160000 ;
      RECT 2.530000 116.080000 4.595000 117.160000 ;
      RECT 1.000000 115.190000 199.100000 116.080000 ;
      RECT 0.000000 114.440000 200.100000 115.190000 ;
      RECT 197.570000 114.340000 200.100000 114.440000 ;
      RECT 0.000000 114.340000 2.530000 114.440000 ;
      RECT 197.570000 113.360000 199.100000 114.340000 ;
      RECT 188.560000 113.360000 195.770000 114.440000 ;
      RECT 143.560000 113.360000 186.760000 114.440000 ;
      RECT 98.560000 113.360000 141.760000 114.440000 ;
      RECT 53.560000 113.360000 96.760000 114.440000 ;
      RECT 8.560000 113.360000 51.760000 114.440000 ;
      RECT 4.330000 113.360000 6.760000 114.440000 ;
      RECT 1.000000 113.360000 2.530000 114.340000 ;
      RECT 0.000000 113.120000 200.100000 113.360000 ;
      RECT 1.000000 112.140000 199.100000 113.120000 ;
      RECT 0.000000 111.720000 200.100000 112.140000 ;
      RECT 199.370000 111.290000 200.100000 111.720000 ;
      RECT 0.000000 111.290000 0.730000 111.720000 ;
      RECT 186.560000 110.640000 197.570000 111.720000 ;
      RECT 141.560000 110.640000 184.760000 111.720000 ;
      RECT 96.560000 110.640000 139.760000 111.720000 ;
      RECT 51.560000 110.640000 94.760000 111.720000 ;
      RECT 6.560000 110.640000 49.760000 111.720000 ;
      RECT 2.530000 110.640000 4.595000 111.720000 ;
      RECT 1.000000 110.310000 199.100000 110.640000 ;
      RECT 0.000000 110.070000 200.100000 110.310000 ;
      RECT 1.000000 109.090000 199.100000 110.070000 ;
      RECT 0.000000 109.000000 200.100000 109.090000 ;
      RECT 197.570000 108.240000 200.100000 109.000000 ;
      RECT 0.000000 108.240000 2.530000 109.000000 ;
      RECT 197.570000 107.920000 199.100000 108.240000 ;
      RECT 188.560000 107.920000 195.770000 109.000000 ;
      RECT 143.560000 107.920000 186.760000 109.000000 ;
      RECT 98.560000 107.920000 141.760000 109.000000 ;
      RECT 53.560000 107.920000 96.760000 109.000000 ;
      RECT 8.560000 107.920000 51.760000 109.000000 ;
      RECT 4.330000 107.920000 6.760000 109.000000 ;
      RECT 1.000000 107.920000 2.530000 108.240000 ;
      RECT 1.000000 107.260000 199.100000 107.920000 ;
      RECT 0.000000 107.020000 200.100000 107.260000 ;
      RECT 1.000000 106.280000 199.100000 107.020000 ;
      RECT 199.370000 105.800000 200.100000 106.040000 ;
      RECT 0.000000 105.800000 0.730000 106.040000 ;
      RECT 186.560000 105.200000 197.570000 106.280000 ;
      RECT 141.560000 105.200000 184.760000 106.280000 ;
      RECT 96.560000 105.200000 139.760000 106.280000 ;
      RECT 51.560000 105.200000 94.760000 106.280000 ;
      RECT 6.560000 105.200000 49.760000 106.280000 ;
      RECT 2.530000 105.200000 4.595000 106.280000 ;
      RECT 1.000000 104.820000 199.100000 105.200000 ;
      RECT 0.000000 103.970000 200.100000 104.820000 ;
      RECT 1.000000 103.560000 199.100000 103.970000 ;
      RECT 197.570000 102.990000 199.100000 103.560000 ;
      RECT 1.000000 102.990000 2.530000 103.560000 ;
      RECT 197.570000 102.750000 200.100000 102.990000 ;
      RECT 0.000000 102.750000 2.530000 102.990000 ;
      RECT 197.570000 102.480000 199.100000 102.750000 ;
      RECT 188.560000 102.480000 195.770000 103.560000 ;
      RECT 143.560000 102.480000 186.760000 103.560000 ;
      RECT 98.560000 102.480000 141.760000 103.560000 ;
      RECT 53.560000 102.480000 96.760000 103.560000 ;
      RECT 8.560000 102.480000 51.760000 103.560000 ;
      RECT 4.330000 102.480000 6.760000 103.560000 ;
      RECT 1.000000 102.480000 2.530000 102.750000 ;
      RECT 1.000000 101.770000 199.100000 102.480000 ;
      RECT 0.000000 100.920000 200.100000 101.770000 ;
      RECT 1.000000 100.840000 199.100000 100.920000 ;
      RECT 199.370000 99.760000 200.100000 99.940000 ;
      RECT 186.560000 99.760000 197.570000 100.840000 ;
      RECT 141.560000 99.760000 184.760000 100.840000 ;
      RECT 96.560000 99.760000 139.760000 100.840000 ;
      RECT 51.560000 99.760000 94.760000 100.840000 ;
      RECT 6.560000 99.760000 49.760000 100.840000 ;
      RECT 2.530000 99.760000 4.595000 100.840000 ;
      RECT 0.000000 99.760000 0.730000 99.940000 ;
      RECT 0.000000 99.700000 200.100000 99.760000 ;
      RECT 1.000000 98.720000 199.100000 99.700000 ;
      RECT 0.000000 98.120000 200.100000 98.720000 ;
      RECT 197.570000 97.870000 200.100000 98.120000 ;
      RECT 0.000000 97.870000 2.530000 98.120000 ;
      RECT 197.570000 97.040000 199.100000 97.870000 ;
      RECT 188.560000 97.040000 195.770000 98.120000 ;
      RECT 143.560000 97.040000 186.760000 98.120000 ;
      RECT 98.560000 97.040000 141.760000 98.120000 ;
      RECT 53.560000 97.040000 96.760000 98.120000 ;
      RECT 8.560000 97.040000 51.760000 98.120000 ;
      RECT 4.330000 97.040000 6.760000 98.120000 ;
      RECT 1.000000 97.040000 2.530000 97.870000 ;
      RECT 1.000000 96.890000 199.100000 97.040000 ;
      RECT 0.000000 96.650000 200.100000 96.890000 ;
      RECT 1.000000 95.670000 199.100000 96.650000 ;
      RECT 0.000000 95.400000 200.100000 95.670000 ;
      RECT 199.370000 94.820000 200.100000 95.400000 ;
      RECT 0.000000 94.820000 0.730000 95.400000 ;
      RECT 186.560000 94.320000 197.570000 95.400000 ;
      RECT 141.560000 94.320000 184.760000 95.400000 ;
      RECT 96.560000 94.320000 139.760000 95.400000 ;
      RECT 51.560000 94.320000 94.760000 95.400000 ;
      RECT 6.560000 94.320000 49.760000 95.400000 ;
      RECT 2.530000 94.320000 4.595000 95.400000 ;
      RECT 1.000000 93.840000 199.100000 94.320000 ;
      RECT 0.000000 93.600000 200.100000 93.840000 ;
      RECT 1.000000 92.680000 199.100000 93.600000 ;
      RECT 197.570000 92.620000 199.100000 92.680000 ;
      RECT 1.000000 92.620000 2.530000 92.680000 ;
      RECT 197.570000 92.380000 200.100000 92.620000 ;
      RECT 0.000000 92.380000 2.530000 92.620000 ;
      RECT 197.570000 91.600000 199.100000 92.380000 ;
      RECT 188.560000 91.600000 195.770000 92.680000 ;
      RECT 143.560000 91.600000 186.760000 92.680000 ;
      RECT 98.560000 91.600000 141.760000 92.680000 ;
      RECT 53.560000 91.600000 96.760000 92.680000 ;
      RECT 8.560000 91.600000 51.760000 92.680000 ;
      RECT 4.330000 91.600000 6.760000 92.680000 ;
      RECT 1.000000 91.600000 2.530000 92.380000 ;
      RECT 1.000000 91.400000 199.100000 91.600000 ;
      RECT 0.000000 90.550000 200.100000 91.400000 ;
      RECT 1.000000 89.960000 199.100000 90.550000 ;
      RECT 199.370000 89.330000 200.100000 89.570000 ;
      RECT 0.000000 89.330000 0.730000 89.570000 ;
      RECT 186.560000 88.880000 197.570000 89.960000 ;
      RECT 141.560000 88.880000 184.760000 89.960000 ;
      RECT 96.560000 88.880000 139.760000 89.960000 ;
      RECT 51.560000 88.880000 94.760000 89.960000 ;
      RECT 6.560000 88.880000 49.760000 89.960000 ;
      RECT 2.530000 88.880000 4.595000 89.960000 ;
      RECT 1.000000 88.350000 199.100000 88.880000 ;
      RECT 0.000000 87.500000 200.100000 88.350000 ;
      RECT 1.000000 87.240000 199.100000 87.500000 ;
      RECT 197.570000 86.520000 199.100000 87.240000 ;
      RECT 1.000000 86.520000 2.530000 87.240000 ;
      RECT 197.570000 86.280000 200.100000 86.520000 ;
      RECT 0.000000 86.280000 2.530000 86.520000 ;
      RECT 197.570000 86.160000 199.100000 86.280000 ;
      RECT 188.560000 86.160000 195.770000 87.240000 ;
      RECT 143.560000 86.160000 186.760000 87.240000 ;
      RECT 98.560000 86.160000 141.760000 87.240000 ;
      RECT 53.560000 86.160000 96.760000 87.240000 ;
      RECT 8.560000 86.160000 51.760000 87.240000 ;
      RECT 4.330000 86.160000 6.760000 87.240000 ;
      RECT 1.000000 86.160000 2.530000 86.280000 ;
      RECT 1.000000 85.300000 199.100000 86.160000 ;
      RECT 0.000000 84.520000 200.100000 85.300000 ;
      RECT 199.370000 84.450000 200.100000 84.520000 ;
      RECT 0.000000 84.450000 0.730000 84.520000 ;
      RECT 199.370000 83.440000 200.100000 83.470000 ;
      RECT 186.560000 83.440000 197.570000 84.520000 ;
      RECT 141.560000 83.440000 184.760000 84.520000 ;
      RECT 96.560000 83.440000 139.760000 84.520000 ;
      RECT 51.560000 83.440000 94.760000 84.520000 ;
      RECT 6.560000 83.440000 49.760000 84.520000 ;
      RECT 2.530000 83.440000 4.595000 84.520000 ;
      RECT 0.000000 83.440000 0.730000 83.470000 ;
      RECT 0.000000 83.230000 200.100000 83.440000 ;
      RECT 1.000000 82.250000 199.100000 83.230000 ;
      RECT 0.000000 81.800000 200.100000 82.250000 ;
      RECT 197.570000 81.400000 200.100000 81.800000 ;
      RECT 0.000000 81.400000 2.530000 81.800000 ;
      RECT 197.570000 80.720000 199.100000 81.400000 ;
      RECT 188.560000 80.720000 195.770000 81.800000 ;
      RECT 143.560000 80.720000 186.760000 81.800000 ;
      RECT 98.560000 80.720000 141.760000 81.800000 ;
      RECT 53.560000 80.720000 96.760000 81.800000 ;
      RECT 8.560000 80.720000 51.760000 81.800000 ;
      RECT 4.330000 80.720000 6.760000 81.800000 ;
      RECT 1.000000 80.720000 2.530000 81.400000 ;
      RECT 1.000000 80.420000 199.100000 80.720000 ;
      RECT 0.000000 80.180000 200.100000 80.420000 ;
      RECT 1.000000 79.200000 199.100000 80.180000 ;
      RECT 0.000000 79.080000 200.100000 79.200000 ;
      RECT 199.370000 78.350000 200.100000 79.080000 ;
      RECT 0.000000 78.350000 0.730000 79.080000 ;
      RECT 186.560000 78.000000 197.570000 79.080000 ;
      RECT 141.560000 78.000000 184.760000 79.080000 ;
      RECT 96.560000 78.000000 139.760000 79.080000 ;
      RECT 51.560000 78.000000 94.760000 79.080000 ;
      RECT 6.560000 78.000000 49.760000 79.080000 ;
      RECT 2.530000 78.000000 4.595000 79.080000 ;
      RECT 1.000000 77.370000 199.100000 78.000000 ;
      RECT 0.000000 77.130000 200.100000 77.370000 ;
      RECT 1.000000 76.360000 199.100000 77.130000 ;
      RECT 197.570000 76.150000 199.100000 76.360000 ;
      RECT 1.000000 76.150000 2.530000 76.360000 ;
      RECT 197.570000 75.910000 200.100000 76.150000 ;
      RECT 0.000000 75.910000 2.530000 76.150000 ;
      RECT 197.570000 75.280000 199.100000 75.910000 ;
      RECT 188.560000 75.280000 195.770000 76.360000 ;
      RECT 143.560000 75.280000 186.760000 76.360000 ;
      RECT 98.560000 75.280000 141.760000 76.360000 ;
      RECT 53.560000 75.280000 96.760000 76.360000 ;
      RECT 8.560000 75.280000 51.760000 76.360000 ;
      RECT 4.330000 75.280000 6.760000 76.360000 ;
      RECT 1.000000 75.280000 2.530000 75.910000 ;
      RECT 1.000000 74.930000 199.100000 75.280000 ;
      RECT 0.000000 74.080000 200.100000 74.930000 ;
      RECT 1.000000 73.640000 199.100000 74.080000 ;
      RECT 199.370000 72.860000 200.100000 73.100000 ;
      RECT 0.000000 72.860000 0.730000 73.100000 ;
      RECT 186.560000 72.560000 197.570000 73.640000 ;
      RECT 141.560000 72.560000 184.760000 73.640000 ;
      RECT 96.560000 72.560000 139.760000 73.640000 ;
      RECT 51.560000 72.560000 94.760000 73.640000 ;
      RECT 6.560000 72.560000 49.760000 73.640000 ;
      RECT 2.530000 72.560000 4.595000 73.640000 ;
      RECT 1.000000 71.880000 199.100000 72.560000 ;
      RECT 0.000000 71.030000 200.100000 71.880000 ;
      RECT 1.000000 70.920000 199.100000 71.030000 ;
      RECT 197.570000 70.050000 199.100000 70.920000 ;
      RECT 1.000000 70.050000 2.530000 70.920000 ;
      RECT 197.570000 69.840000 200.100000 70.050000 ;
      RECT 188.560000 69.840000 195.770000 70.920000 ;
      RECT 143.560000 69.840000 186.760000 70.920000 ;
      RECT 98.560000 69.840000 141.760000 70.920000 ;
      RECT 53.560000 69.840000 96.760000 70.920000 ;
      RECT 8.560000 69.840000 51.760000 70.920000 ;
      RECT 4.330000 69.840000 6.760000 70.920000 ;
      RECT 0.000000 69.840000 2.530000 70.050000 ;
      RECT 0.000000 69.810000 200.100000 69.840000 ;
      RECT 1.000000 68.830000 199.100000 69.810000 ;
      RECT 0.000000 68.200000 200.100000 68.830000 ;
      RECT 199.370000 67.980000 200.100000 68.200000 ;
      RECT 0.000000 67.980000 0.730000 68.200000 ;
      RECT 186.560000 67.120000 197.570000 68.200000 ;
      RECT 141.560000 67.120000 184.760000 68.200000 ;
      RECT 96.560000 67.120000 139.760000 68.200000 ;
      RECT 51.560000 67.120000 94.760000 68.200000 ;
      RECT 6.560000 67.120000 49.760000 68.200000 ;
      RECT 2.530000 67.120000 4.595000 68.200000 ;
      RECT 1.000000 67.000000 199.100000 67.120000 ;
      RECT 0.000000 66.760000 200.100000 67.000000 ;
      RECT 1.000000 65.780000 199.100000 66.760000 ;
      RECT 0.000000 65.480000 200.100000 65.780000 ;
      RECT 197.570000 64.930000 200.100000 65.480000 ;
      RECT 0.000000 64.930000 2.530000 65.480000 ;
      RECT 197.570000 64.400000 199.100000 64.930000 ;
      RECT 188.560000 64.400000 195.770000 65.480000 ;
      RECT 143.560000 64.400000 186.760000 65.480000 ;
      RECT 98.560000 64.400000 141.760000 65.480000 ;
      RECT 53.560000 64.400000 96.760000 65.480000 ;
      RECT 8.560000 64.400000 51.760000 65.480000 ;
      RECT 4.330000 64.400000 6.760000 65.480000 ;
      RECT 1.000000 64.400000 2.530000 64.930000 ;
      RECT 1.000000 63.950000 199.100000 64.400000 ;
      RECT 0.000000 63.710000 200.100000 63.950000 ;
      RECT 1.000000 62.760000 199.100000 63.710000 ;
      RECT 199.370000 62.490000 200.100000 62.730000 ;
      RECT 0.000000 62.490000 0.730000 62.730000 ;
      RECT 186.560000 61.680000 197.570000 62.760000 ;
      RECT 141.560000 61.680000 184.760000 62.760000 ;
      RECT 96.560000 61.680000 139.760000 62.760000 ;
      RECT 51.560000 61.680000 94.760000 62.760000 ;
      RECT 6.560000 61.680000 49.760000 62.760000 ;
      RECT 2.530000 61.680000 4.595000 62.760000 ;
      RECT 1.000000 61.510000 199.100000 61.680000 ;
      RECT 0.000000 60.660000 200.100000 61.510000 ;
      RECT 1.000000 60.040000 199.100000 60.660000 ;
      RECT 197.570000 59.680000 199.100000 60.040000 ;
      RECT 1.000000 59.680000 2.530000 60.040000 ;
      RECT 197.570000 59.440000 200.100000 59.680000 ;
      RECT 0.000000 59.440000 2.530000 59.680000 ;
      RECT 197.570000 58.960000 199.100000 59.440000 ;
      RECT 188.560000 58.960000 195.770000 60.040000 ;
      RECT 143.560000 58.960000 186.760000 60.040000 ;
      RECT 98.560000 58.960000 141.760000 60.040000 ;
      RECT 53.560000 58.960000 96.760000 60.040000 ;
      RECT 8.560000 58.960000 51.760000 60.040000 ;
      RECT 4.330000 58.960000 6.760000 60.040000 ;
      RECT 1.000000 58.960000 2.530000 59.440000 ;
      RECT 1.000000 58.460000 199.100000 58.960000 ;
      RECT 0.000000 57.610000 200.100000 58.460000 ;
      RECT 1.000000 57.320000 199.100000 57.610000 ;
      RECT 199.370000 56.390000 200.100000 56.630000 ;
      RECT 0.000000 56.390000 0.730000 56.630000 ;
      RECT 186.560000 56.240000 197.570000 57.320000 ;
      RECT 141.560000 56.240000 184.760000 57.320000 ;
      RECT 96.560000 56.240000 139.760000 57.320000 ;
      RECT 51.560000 56.240000 94.760000 57.320000 ;
      RECT 6.560000 56.240000 49.760000 57.320000 ;
      RECT 2.530000 56.240000 4.595000 57.320000 ;
      RECT 1.000000 55.410000 199.100000 56.240000 ;
      RECT 0.000000 54.600000 200.100000 55.410000 ;
      RECT 197.570000 54.560000 200.100000 54.600000 ;
      RECT 0.000000 54.560000 2.530000 54.600000 ;
      RECT 197.570000 53.580000 199.100000 54.560000 ;
      RECT 1.000000 53.580000 2.530000 54.560000 ;
      RECT 197.570000 53.520000 200.100000 53.580000 ;
      RECT 188.560000 53.520000 195.770000 54.600000 ;
      RECT 143.560000 53.520000 186.760000 54.600000 ;
      RECT 98.560000 53.520000 141.760000 54.600000 ;
      RECT 53.560000 53.520000 96.760000 54.600000 ;
      RECT 8.560000 53.520000 51.760000 54.600000 ;
      RECT 4.330000 53.520000 6.760000 54.600000 ;
      RECT 0.000000 53.520000 2.530000 53.580000 ;
      RECT 0.000000 53.340000 200.100000 53.520000 ;
      RECT 1.000000 52.360000 199.100000 53.340000 ;
      RECT 0.000000 51.880000 200.100000 52.360000 ;
      RECT 199.370000 51.510000 200.100000 51.880000 ;
      RECT 0.000000 51.510000 0.730000 51.880000 ;
      RECT 186.560000 50.800000 197.570000 51.880000 ;
      RECT 141.560000 50.800000 184.760000 51.880000 ;
      RECT 96.560000 50.800000 139.760000 51.880000 ;
      RECT 51.560000 50.800000 94.760000 51.880000 ;
      RECT 6.560000 50.800000 49.760000 51.880000 ;
      RECT 2.530000 50.800000 4.595000 51.880000 ;
      RECT 1.000000 50.530000 199.100000 50.800000 ;
      RECT 0.000000 50.290000 200.100000 50.530000 ;
      RECT 1.000000 49.310000 199.100000 50.290000 ;
      RECT 0.000000 49.160000 200.100000 49.310000 ;
      RECT 197.570000 49.070000 200.100000 49.160000 ;
      RECT 0.000000 49.070000 2.530000 49.160000 ;
      RECT 197.570000 48.090000 199.100000 49.070000 ;
      RECT 1.000000 48.090000 2.530000 49.070000 ;
      RECT 197.570000 48.080000 200.100000 48.090000 ;
      RECT 188.560000 48.080000 195.770000 49.160000 ;
      RECT 143.560000 48.080000 186.760000 49.160000 ;
      RECT 98.560000 48.080000 141.760000 49.160000 ;
      RECT 53.560000 48.080000 96.760000 49.160000 ;
      RECT 8.560000 48.080000 51.760000 49.160000 ;
      RECT 4.330000 48.080000 6.760000 49.160000 ;
      RECT 0.000000 48.080000 2.530000 48.090000 ;
      RECT 0.000000 47.240000 200.100000 48.080000 ;
      RECT 1.000000 46.440000 199.100000 47.240000 ;
      RECT 199.370000 46.020000 200.100000 46.260000 ;
      RECT 0.000000 46.020000 0.730000 46.260000 ;
      RECT 186.560000 45.360000 197.570000 46.440000 ;
      RECT 141.560000 45.360000 184.760000 46.440000 ;
      RECT 96.560000 45.360000 139.760000 46.440000 ;
      RECT 51.560000 45.360000 94.760000 46.440000 ;
      RECT 6.560000 45.360000 49.760000 46.440000 ;
      RECT 2.530000 45.360000 4.595000 46.440000 ;
      RECT 1.000000 45.040000 199.100000 45.360000 ;
      RECT 0.000000 44.190000 200.100000 45.040000 ;
      RECT 1.000000 43.720000 199.100000 44.190000 ;
      RECT 197.570000 43.210000 199.100000 43.720000 ;
      RECT 1.000000 43.210000 2.530000 43.720000 ;
      RECT 197.570000 42.970000 200.100000 43.210000 ;
      RECT 0.000000 42.970000 2.530000 43.210000 ;
      RECT 197.570000 42.640000 199.100000 42.970000 ;
      RECT 188.560000 42.640000 195.770000 43.720000 ;
      RECT 143.560000 42.640000 186.760000 43.720000 ;
      RECT 98.560000 42.640000 141.760000 43.720000 ;
      RECT 53.560000 42.640000 96.760000 43.720000 ;
      RECT 8.560000 42.640000 51.760000 43.720000 ;
      RECT 4.330000 42.640000 6.760000 43.720000 ;
      RECT 1.000000 42.640000 2.530000 42.970000 ;
      RECT 1.000000 41.990000 199.100000 42.640000 ;
      RECT 0.000000 41.140000 200.100000 41.990000 ;
      RECT 1.000000 41.000000 199.100000 41.140000 ;
      RECT 199.370000 39.920000 200.100000 40.160000 ;
      RECT 186.560000 39.920000 197.570000 41.000000 ;
      RECT 141.560000 39.920000 184.760000 41.000000 ;
      RECT 96.560000 39.920000 139.760000 41.000000 ;
      RECT 51.560000 39.920000 94.760000 41.000000 ;
      RECT 6.560000 39.920000 49.760000 41.000000 ;
      RECT 2.530000 39.920000 4.595000 41.000000 ;
      RECT 0.000000 39.920000 0.730000 40.160000 ;
      RECT 1.000000 38.940000 199.100000 39.920000 ;
      RECT 0.000000 38.280000 200.100000 38.940000 ;
      RECT 197.570000 38.090000 200.100000 38.280000 ;
      RECT 0.000000 38.090000 2.530000 38.280000 ;
      RECT 197.570000 37.200000 199.100000 38.090000 ;
      RECT 188.560000 37.200000 195.770000 38.280000 ;
      RECT 143.560000 37.200000 186.760000 38.280000 ;
      RECT 98.560000 37.200000 141.760000 38.280000 ;
      RECT 53.560000 37.200000 96.760000 38.280000 ;
      RECT 8.560000 37.200000 51.760000 38.280000 ;
      RECT 4.330000 37.200000 6.760000 38.280000 ;
      RECT 1.000000 37.200000 2.530000 38.090000 ;
      RECT 1.000000 37.110000 199.100000 37.200000 ;
      RECT 0.000000 36.870000 200.100000 37.110000 ;
      RECT 1.000000 35.890000 199.100000 36.870000 ;
      RECT 0.000000 35.560000 200.100000 35.890000 ;
      RECT 199.370000 35.040000 200.100000 35.560000 ;
      RECT 0.000000 35.040000 0.730000 35.560000 ;
      RECT 186.560000 34.480000 197.570000 35.560000 ;
      RECT 141.560000 34.480000 184.760000 35.560000 ;
      RECT 96.560000 34.480000 139.760000 35.560000 ;
      RECT 51.560000 34.480000 94.760000 35.560000 ;
      RECT 6.560000 34.480000 49.760000 35.560000 ;
      RECT 2.530000 34.480000 4.595000 35.560000 ;
      RECT 1.000000 34.060000 199.100000 34.480000 ;
      RECT 0.000000 33.820000 200.100000 34.060000 ;
      RECT 1.000000 32.840000 199.100000 33.820000 ;
      RECT 197.570000 32.600000 200.100000 32.840000 ;
      RECT 0.000000 32.600000 2.530000 32.840000 ;
      RECT 197.570000 31.760000 199.100000 32.600000 ;
      RECT 188.560000 31.760000 195.770000 32.840000 ;
      RECT 143.560000 31.760000 186.760000 32.840000 ;
      RECT 98.560000 31.760000 141.760000 32.840000 ;
      RECT 53.560000 31.760000 96.760000 32.840000 ;
      RECT 8.560000 31.760000 51.760000 32.840000 ;
      RECT 4.330000 31.760000 6.760000 32.840000 ;
      RECT 1.000000 31.760000 2.530000 32.600000 ;
      RECT 1.000000 31.620000 199.100000 31.760000 ;
      RECT 0.000000 30.770000 200.100000 31.620000 ;
      RECT 1.000000 30.120000 199.100000 30.770000 ;
      RECT 199.370000 29.550000 200.100000 29.790000 ;
      RECT 0.000000 29.550000 0.730000 29.790000 ;
      RECT 186.560000 29.040000 197.570000 30.120000 ;
      RECT 141.560000 29.040000 184.760000 30.120000 ;
      RECT 96.560000 29.040000 139.760000 30.120000 ;
      RECT 51.560000 29.040000 94.760000 30.120000 ;
      RECT 6.560000 29.040000 49.760000 30.120000 ;
      RECT 2.530000 29.040000 4.595000 30.120000 ;
      RECT 1.000000 28.570000 199.100000 29.040000 ;
      RECT 0.000000 27.720000 200.100000 28.570000 ;
      RECT 1.000000 27.400000 199.100000 27.720000 ;
      RECT 197.570000 26.740000 199.100000 27.400000 ;
      RECT 1.000000 26.740000 2.530000 27.400000 ;
      RECT 197.570000 26.500000 200.100000 26.740000 ;
      RECT 0.000000 26.500000 2.530000 26.740000 ;
      RECT 197.570000 26.320000 199.100000 26.500000 ;
      RECT 188.560000 26.320000 195.770000 27.400000 ;
      RECT 143.560000 26.320000 186.760000 27.400000 ;
      RECT 98.560000 26.320000 141.760000 27.400000 ;
      RECT 53.560000 26.320000 96.760000 27.400000 ;
      RECT 8.560000 26.320000 51.760000 27.400000 ;
      RECT 4.330000 26.320000 6.760000 27.400000 ;
      RECT 1.000000 26.320000 2.530000 26.500000 ;
      RECT 1.000000 25.520000 199.100000 26.320000 ;
      RECT 0.000000 24.680000 200.100000 25.520000 ;
      RECT 199.370000 24.670000 200.100000 24.680000 ;
      RECT 0.000000 24.670000 0.730000 24.680000 ;
      RECT 199.370000 23.600000 200.100000 23.690000 ;
      RECT 186.560000 23.600000 197.570000 24.680000 ;
      RECT 141.560000 23.600000 184.760000 24.680000 ;
      RECT 96.560000 23.600000 139.760000 24.680000 ;
      RECT 51.560000 23.600000 94.760000 24.680000 ;
      RECT 6.560000 23.600000 49.760000 24.680000 ;
      RECT 2.530000 23.600000 4.595000 24.680000 ;
      RECT 0.000000 23.600000 0.730000 23.690000 ;
      RECT 0.000000 23.450000 200.100000 23.600000 ;
      RECT 1.000000 22.470000 199.100000 23.450000 ;
      RECT 0.000000 21.960000 200.100000 22.470000 ;
      RECT 197.570000 21.620000 200.100000 21.960000 ;
      RECT 0.000000 21.620000 2.530000 21.960000 ;
      RECT 197.570000 20.880000 199.100000 21.620000 ;
      RECT 188.560000 20.880000 195.770000 21.960000 ;
      RECT 143.560000 20.880000 186.760000 21.960000 ;
      RECT 98.560000 20.880000 141.760000 21.960000 ;
      RECT 53.560000 20.880000 96.760000 21.960000 ;
      RECT 8.560000 20.880000 51.760000 21.960000 ;
      RECT 4.330000 20.880000 6.760000 21.960000 ;
      RECT 1.000000 20.880000 2.530000 21.620000 ;
      RECT 1.000000 20.640000 199.100000 20.880000 ;
      RECT 0.000000 20.400000 200.100000 20.640000 ;
      RECT 1.000000 19.420000 199.100000 20.400000 ;
      RECT 0.000000 19.240000 200.100000 19.420000 ;
      RECT 199.370000 19.180000 200.100000 19.240000 ;
      RECT 0.000000 19.180000 0.730000 19.240000 ;
      RECT 199.370000 18.160000 200.100000 18.200000 ;
      RECT 186.560000 18.160000 197.570000 19.240000 ;
      RECT 141.560000 18.160000 184.760000 19.240000 ;
      RECT 96.560000 18.160000 139.760000 19.240000 ;
      RECT 51.560000 18.160000 94.760000 19.240000 ;
      RECT 6.560000 18.160000 49.760000 19.240000 ;
      RECT 2.530000 18.160000 4.595000 19.240000 ;
      RECT 0.000000 18.160000 0.730000 18.200000 ;
      RECT 0.000000 17.350000 200.100000 18.160000 ;
      RECT 1.000000 16.520000 199.100000 17.350000 ;
      RECT 197.570000 16.370000 199.100000 16.520000 ;
      RECT 1.000000 16.370000 2.530000 16.520000 ;
      RECT 197.570000 16.130000 200.100000 16.370000 ;
      RECT 0.000000 16.130000 2.530000 16.370000 ;
      RECT 197.570000 15.440000 199.100000 16.130000 ;
      RECT 188.560000 15.440000 195.770000 16.520000 ;
      RECT 143.560000 15.440000 186.760000 16.520000 ;
      RECT 98.560000 15.440000 141.760000 16.520000 ;
      RECT 53.560000 15.440000 96.760000 16.520000 ;
      RECT 8.560000 15.440000 51.760000 16.520000 ;
      RECT 4.330000 15.440000 6.760000 16.520000 ;
      RECT 1.000000 15.440000 2.530000 16.130000 ;
      RECT 1.000000 15.150000 199.100000 15.440000 ;
      RECT 0.000000 14.300000 200.100000 15.150000 ;
      RECT 1.000000 13.800000 199.100000 14.300000 ;
      RECT 199.370000 13.080000 200.100000 13.320000 ;
      RECT 0.000000 13.080000 0.730000 13.320000 ;
      RECT 186.560000 12.720000 197.570000 13.800000 ;
      RECT 141.560000 12.720000 184.760000 13.800000 ;
      RECT 96.560000 12.720000 139.760000 13.800000 ;
      RECT 51.560000 12.720000 94.760000 13.800000 ;
      RECT 6.560000 12.720000 49.760000 13.800000 ;
      RECT 2.530000 12.720000 4.595000 13.800000 ;
      RECT 1.000000 12.100000 199.100000 12.720000 ;
      RECT 0.000000 11.250000 200.100000 12.100000 ;
      RECT 1.000000 11.080000 199.100000 11.250000 ;
      RECT 197.570000 10.270000 199.100000 11.080000 ;
      RECT 1.000000 10.270000 2.530000 11.080000 ;
      RECT 197.570000 10.030000 200.100000 10.270000 ;
      RECT 0.000000 10.030000 2.530000 10.270000 ;
      RECT 197.570000 10.000000 199.100000 10.030000 ;
      RECT 188.560000 10.000000 195.770000 11.080000 ;
      RECT 143.560000 10.000000 186.760000 11.080000 ;
      RECT 98.560000 10.000000 141.760000 11.080000 ;
      RECT 53.560000 10.000000 96.760000 11.080000 ;
      RECT 8.560000 10.000000 51.760000 11.080000 ;
      RECT 4.330000 10.000000 6.760000 11.080000 ;
      RECT 1.000000 10.000000 2.530000 10.030000 ;
      RECT 1.000000 9.050000 199.100000 10.000000 ;
      RECT 0.000000 8.360000 200.100000 9.050000 ;
      RECT 199.370000 8.200000 200.100000 8.360000 ;
      RECT 0.000000 8.200000 0.730000 8.360000 ;
      RECT 186.560000 7.280000 197.570000 8.360000 ;
      RECT 141.560000 7.280000 184.760000 8.360000 ;
      RECT 96.560000 7.280000 139.760000 8.360000 ;
      RECT 51.560000 7.280000 94.760000 8.360000 ;
      RECT 6.560000 7.280000 49.760000 8.360000 ;
      RECT 2.530000 7.280000 4.595000 8.360000 ;
      RECT 1.000000 7.220000 199.100000 7.280000 ;
      RECT 0.000000 6.980000 200.100000 7.220000 ;
      RECT 1.000000 6.000000 199.100000 6.980000 ;
      RECT 0.000000 5.760000 200.100000 6.000000 ;
      RECT 1.000000 5.640000 199.100000 5.760000 ;
      RECT 197.570000 4.780000 199.100000 5.640000 ;
      RECT 1.000000 4.780000 2.530000 5.640000 ;
      RECT 197.570000 4.560000 200.100000 4.780000 ;
      RECT 188.560000 4.560000 195.770000 5.640000 ;
      RECT 143.560000 4.560000 186.760000 5.640000 ;
      RECT 98.560000 4.560000 141.760000 5.640000 ;
      RECT 53.560000 4.560000 96.760000 5.640000 ;
      RECT 8.560000 4.560000 51.760000 5.640000 ;
      RECT 4.330000 4.560000 6.760000 5.640000 ;
      RECT 0.000000 4.560000 2.530000 4.780000 ;
      RECT 0.000000 4.350000 200.100000 4.560000 ;
      RECT 0.000000 0.000000 200.100000 0.750000 ;
    LAYER met4 ;
      RECT 4.330000 399.090000 195.770000 400.520000 ;
      RECT 186.560000 397.290000 195.770000 399.090000 ;
      RECT 141.560000 397.290000 184.760000 399.090000 ;
      RECT 96.560000 397.290000 139.760000 399.090000 ;
      RECT 51.560000 397.290000 94.760000 399.090000 ;
      RECT 6.560000 397.290000 49.760000 399.090000 ;
      RECT 4.330000 394.600000 4.760000 399.090000 ;
      RECT 4.330000 393.520000 4.595000 394.600000 ;
      RECT 4.330000 389.160000 4.760000 393.520000 ;
      RECT 4.330000 388.080000 4.595000 389.160000 ;
      RECT 4.330000 383.720000 4.760000 388.080000 ;
      RECT 4.330000 382.640000 4.595000 383.720000 ;
      RECT 4.330000 378.280000 4.760000 382.640000 ;
      RECT 4.330000 377.200000 4.595000 378.280000 ;
      RECT 4.330000 372.840000 4.760000 377.200000 ;
      RECT 4.330000 371.760000 4.595000 372.840000 ;
      RECT 4.330000 367.400000 4.760000 371.760000 ;
      RECT 4.330000 366.320000 4.595000 367.400000 ;
      RECT 4.330000 361.960000 4.760000 366.320000 ;
      RECT 4.330000 360.880000 4.595000 361.960000 ;
      RECT 4.330000 356.520000 4.760000 360.880000 ;
      RECT 4.330000 355.440000 4.595000 356.520000 ;
      RECT 4.330000 351.080000 4.760000 355.440000 ;
      RECT 4.330000 350.000000 4.595000 351.080000 ;
      RECT 4.330000 345.640000 4.760000 350.000000 ;
      RECT 4.330000 344.560000 4.595000 345.640000 ;
      RECT 4.330000 340.200000 4.760000 344.560000 ;
      RECT 4.330000 339.120000 4.595000 340.200000 ;
      RECT 4.330000 334.760000 4.760000 339.120000 ;
      RECT 4.330000 333.680000 4.595000 334.760000 ;
      RECT 4.330000 329.320000 4.760000 333.680000 ;
      RECT 4.330000 328.240000 4.595000 329.320000 ;
      RECT 4.330000 323.880000 4.760000 328.240000 ;
      RECT 4.330000 322.800000 4.595000 323.880000 ;
      RECT 4.330000 318.440000 4.760000 322.800000 ;
      RECT 4.330000 317.360000 4.595000 318.440000 ;
      RECT 4.330000 313.000000 4.760000 317.360000 ;
      RECT 4.330000 311.920000 4.595000 313.000000 ;
      RECT 4.330000 307.560000 4.760000 311.920000 ;
      RECT 4.330000 306.480000 4.595000 307.560000 ;
      RECT 4.330000 302.120000 4.760000 306.480000 ;
      RECT 4.330000 301.040000 4.595000 302.120000 ;
      RECT 4.330000 296.680000 4.760000 301.040000 ;
      RECT 4.330000 295.600000 4.595000 296.680000 ;
      RECT 4.330000 291.240000 4.760000 295.600000 ;
      RECT 4.330000 290.160000 4.595000 291.240000 ;
      RECT 4.330000 285.800000 4.760000 290.160000 ;
      RECT 4.330000 284.720000 4.595000 285.800000 ;
      RECT 4.330000 280.360000 4.760000 284.720000 ;
      RECT 4.330000 279.280000 4.595000 280.360000 ;
      RECT 4.330000 274.920000 4.760000 279.280000 ;
      RECT 4.330000 273.840000 4.595000 274.920000 ;
      RECT 4.330000 269.480000 4.760000 273.840000 ;
      RECT 4.330000 268.400000 4.595000 269.480000 ;
      RECT 4.330000 264.040000 4.760000 268.400000 ;
      RECT 4.330000 262.960000 4.595000 264.040000 ;
      RECT 4.330000 258.600000 4.760000 262.960000 ;
      RECT 4.330000 257.520000 4.595000 258.600000 ;
      RECT 4.330000 253.160000 4.760000 257.520000 ;
      RECT 4.330000 252.080000 4.595000 253.160000 ;
      RECT 4.330000 247.720000 4.760000 252.080000 ;
      RECT 4.330000 246.640000 4.595000 247.720000 ;
      RECT 4.330000 242.280000 4.760000 246.640000 ;
      RECT 4.330000 241.200000 4.595000 242.280000 ;
      RECT 4.330000 236.840000 4.760000 241.200000 ;
      RECT 4.330000 235.760000 4.595000 236.840000 ;
      RECT 4.330000 231.400000 4.760000 235.760000 ;
      RECT 4.330000 230.320000 4.595000 231.400000 ;
      RECT 4.330000 225.960000 4.760000 230.320000 ;
      RECT 4.330000 224.880000 4.595000 225.960000 ;
      RECT 4.330000 220.520000 4.760000 224.880000 ;
      RECT 4.330000 219.440000 4.595000 220.520000 ;
      RECT 4.330000 215.080000 4.760000 219.440000 ;
      RECT 4.330000 214.000000 4.595000 215.080000 ;
      RECT 4.330000 209.640000 4.760000 214.000000 ;
      RECT 4.330000 208.560000 4.595000 209.640000 ;
      RECT 4.330000 204.200000 4.760000 208.560000 ;
      RECT 4.330000 203.120000 4.595000 204.200000 ;
      RECT 4.330000 198.760000 4.760000 203.120000 ;
      RECT 4.330000 197.680000 4.595000 198.760000 ;
      RECT 4.330000 193.320000 4.760000 197.680000 ;
      RECT 4.330000 192.240000 4.595000 193.320000 ;
      RECT 4.330000 187.880000 4.760000 192.240000 ;
      RECT 4.330000 186.800000 4.595000 187.880000 ;
      RECT 4.330000 182.440000 4.760000 186.800000 ;
      RECT 4.330000 181.360000 4.595000 182.440000 ;
      RECT 4.330000 177.000000 4.760000 181.360000 ;
      RECT 4.330000 175.920000 4.595000 177.000000 ;
      RECT 4.330000 171.560000 4.760000 175.920000 ;
      RECT 4.330000 170.480000 4.595000 171.560000 ;
      RECT 4.330000 166.120000 4.760000 170.480000 ;
      RECT 4.330000 165.040000 4.595000 166.120000 ;
      RECT 4.330000 160.680000 4.760000 165.040000 ;
      RECT 4.330000 159.600000 4.595000 160.680000 ;
      RECT 4.330000 155.240000 4.760000 159.600000 ;
      RECT 4.330000 154.160000 4.595000 155.240000 ;
      RECT 4.330000 149.800000 4.760000 154.160000 ;
      RECT 4.330000 148.720000 4.595000 149.800000 ;
      RECT 4.330000 144.360000 4.760000 148.720000 ;
      RECT 4.330000 143.280000 4.595000 144.360000 ;
      RECT 4.330000 138.920000 4.760000 143.280000 ;
      RECT 4.330000 137.840000 4.595000 138.920000 ;
      RECT 4.330000 133.480000 4.760000 137.840000 ;
      RECT 4.330000 132.400000 4.595000 133.480000 ;
      RECT 4.330000 128.040000 4.760000 132.400000 ;
      RECT 4.330000 126.960000 4.595000 128.040000 ;
      RECT 4.330000 122.600000 4.760000 126.960000 ;
      RECT 4.330000 121.520000 4.595000 122.600000 ;
      RECT 4.330000 117.160000 4.760000 121.520000 ;
      RECT 4.330000 116.080000 4.595000 117.160000 ;
      RECT 4.330000 111.720000 4.760000 116.080000 ;
      RECT 4.330000 110.640000 4.595000 111.720000 ;
      RECT 4.330000 106.280000 4.760000 110.640000 ;
      RECT 4.330000 105.200000 4.595000 106.280000 ;
      RECT 4.330000 100.840000 4.760000 105.200000 ;
      RECT 4.330000 99.760000 4.595000 100.840000 ;
      RECT 4.330000 95.400000 4.760000 99.760000 ;
      RECT 4.330000 94.320000 4.595000 95.400000 ;
      RECT 4.330000 89.960000 4.760000 94.320000 ;
      RECT 4.330000 88.880000 4.595000 89.960000 ;
      RECT 4.330000 84.520000 4.760000 88.880000 ;
      RECT 4.330000 83.440000 4.595000 84.520000 ;
      RECT 4.330000 79.080000 4.760000 83.440000 ;
      RECT 4.330000 78.000000 4.595000 79.080000 ;
      RECT 4.330000 73.640000 4.760000 78.000000 ;
      RECT 4.330000 72.560000 4.595000 73.640000 ;
      RECT 4.330000 68.200000 4.760000 72.560000 ;
      RECT 4.330000 67.120000 4.595000 68.200000 ;
      RECT 4.330000 62.760000 4.760000 67.120000 ;
      RECT 4.330000 61.680000 4.595000 62.760000 ;
      RECT 4.330000 57.320000 4.760000 61.680000 ;
      RECT 4.330000 56.240000 4.595000 57.320000 ;
      RECT 4.330000 51.880000 4.760000 56.240000 ;
      RECT 4.330000 50.800000 4.595000 51.880000 ;
      RECT 4.330000 46.440000 4.760000 50.800000 ;
      RECT 4.330000 45.360000 4.595000 46.440000 ;
      RECT 4.330000 41.000000 4.760000 45.360000 ;
      RECT 4.330000 39.920000 4.595000 41.000000 ;
      RECT 4.330000 35.560000 4.760000 39.920000 ;
      RECT 4.330000 34.480000 4.595000 35.560000 ;
      RECT 4.330000 30.120000 4.760000 34.480000 ;
      RECT 4.330000 29.040000 4.595000 30.120000 ;
      RECT 4.330000 24.680000 4.760000 29.040000 ;
      RECT 4.330000 23.600000 4.595000 24.680000 ;
      RECT 4.330000 19.240000 4.760000 23.600000 ;
      RECT 4.330000 18.160000 4.595000 19.240000 ;
      RECT 4.330000 13.800000 4.760000 18.160000 ;
      RECT 4.330000 12.720000 4.595000 13.800000 ;
      RECT 4.330000 8.360000 4.760000 12.720000 ;
      RECT 4.330000 7.280000 4.595000 8.360000 ;
      RECT 188.560000 2.550000 195.770000 397.290000 ;
      RECT 186.560000 2.550000 186.760000 397.290000 ;
      RECT 143.560000 2.550000 184.760000 397.290000 ;
      RECT 141.560000 2.550000 141.760000 397.290000 ;
      RECT 98.560000 2.550000 139.760000 397.290000 ;
      RECT 96.560000 2.550000 96.760000 397.290000 ;
      RECT 53.560000 2.550000 94.760000 397.290000 ;
      RECT 51.560000 2.550000 51.760000 397.290000 ;
      RECT 8.560000 2.550000 49.760000 397.290000 ;
      RECT 6.560000 2.550000 6.760000 397.290000 ;
      RECT 186.560000 0.750000 195.770000 2.550000 ;
      RECT 141.560000 0.750000 184.760000 2.550000 ;
      RECT 96.560000 0.750000 139.760000 2.550000 ;
      RECT 51.560000 0.750000 94.760000 2.550000 ;
      RECT 6.560000 0.750000 49.760000 2.550000 ;
      RECT 4.330000 0.750000 4.760000 7.280000 ;
      RECT 199.370000 0.000000 200.100000 400.520000 ;
      RECT 4.330000 0.000000 195.770000 0.750000 ;
      RECT 0.000000 0.000000 0.730000 400.520000 ;
  END
END DSP

END LIBRARY
